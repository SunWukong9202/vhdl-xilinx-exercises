----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:10:30 11/21/2022 
-- Design Name: 
-- Module Name:    pong_TOP - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity pong_TOP is
	port(
		i_clk: in std_logic;
		o_R0,o_R1,o_R2: out std_logic;	--RED COLOR	
		o_G0,o_G1,o_G2: out std_logic;	--GREEN COLOR	
		o_B0,o_B1: out std_logic;		--BLUE COLOR
		o_HS: out std_logic;
		o_VS: out std_logic;
		i_joystick_p1: in std_logic_vector(5 downto 0);		
		i_joystick_p2: in std_logic_vector(5 downto 0);
		o_paddle_sound_collide: out std_logic;
		i_select: in std_logic;
		i_difficulty: in std_logic_vector(1 downto 0)
	);
end pong_TOP;

architecture Behavioral of pong_TOP is
	type rom_bitmap is array (0 to 2951) of integer;
	type rom_bitmap_arrow is array (0 to 647) of integer;	
	type rom_bitmap_title is array (0 to 8999) of integer;		
	type rom_bitmap_title_2 is array (0 to 8909) of integer;	
	type rom_bitmap_ball is array (0 to 399) of integer;
	
	constant rom_pong: rom_bitmap_title_2 := (
	0 => 0, 1 => 1, 2 => 1, 3 => 1, 4 => 1, 5 => 1, 6 => 1, 7 => 1, 8 => 1, 9 => 1, 10 => 1, 11 => 1, 12 => 1, 13 => 1, 14 => 1, 15 => 1, 16 => 1, 17 => 1, 18 => 1, 19 => 1, 20 => 1, 21 => 1, 22 => 1, 23 => 1, 24 => 1, 25 => 1, 26 => 1, 27 => 1, 28 => 1, 29 => 1, 30 => 1, 31 => 1, 32 => 1, 33 => 1, 34 => 
1, 35 => 1, 36 => 1, 37 => 0, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 0, 45 => 0, 46 => 0, 47 => 0, 48 => 0, 49 => 0, 50 => 0, 51 => 0, 52 => 0, 53 => 0, 54 => 0, 55 => 0, 56 => 0, 57 => 0, 58 => 1, 59 => 1, 60 => 1, 61 => 1, 62 => 1, 63 => 1, 64 => 1, 65 => 1, 66 => 1, 67 => 1, 68 => 1, 69 => 1, 70 => 1, 71 => 1, 72 => 1, 73 => 1, 74 => 1, 75 => 1, 76 => 1, 77 => 1, 78 => 1, 79 => 1, 80 => 1, 81 => 1, 82 => 1, 83 => 1, 84 => 1, 
85 => 1, 86 => 1, 87 => 1, 88 => 1, 89 => 0, 90 => 0, 91 => 0, 92 => 0, 93 => 0, 94 => 0, 95 => 0, 96 => 0, 97 => 0, 98 => 0, 99 => 0, 100 => 0, 101 => 0, 102 => 0, 103 => 1, 104 => 1, 105 => 1, 106 => 1, 107 => 1, 108 => 0, 109 => 0, 110 => 0, 111 => 0, 112 => 0, 113 => 0, 114 => 0, 115 => 0, 116 => 
0, 117 => 0, 118 => 0, 119 => 0, 120 => 0, 121 => 0, 122 => 0, 123 => 0, 124 => 0, 125 => 0, 126 => 0, 127 => 0, 128 => 0, 129 => 0, 130 => 0, 131 => 0, 132 => 0, 133 => 0, 134 => 0, 135 => 1, 136 => 1, 137 => 1, 138 => 1, 139 => 1, 140 => 1, 141 => 1, 142 => 1, 143 => 1, 144 => 1, 145 => 1, 146 => 0, 147 => 0, 148 => 0, 149 => 0, 150 => 0, 151 => 0, 152 => 0, 153 => 0, 154 => 0, 155 => 0, 156 => 0, 157 => 0, 158 => 0, 159 => 0, 160 => 0, 161 => 1, 
162 => 1, 163 => 1, 164 => 1, 165 => 1, 166 => 1, 167 => 1, 168 => 1, 169 => 1, 170 => 1, 171 => 1, 172 => 1, 173 => 1, 174 => 1, 175 => 1, 176 => 1, 177 => 1, 178 => 1, 179 => 1, 180 => 1, 181 => 1, 182 => 1, 183 => 1, 184 => 1, 185 => 1, 186 => 1, 187 => 1, 188 => 1, 189 => 1, 190 => 1, 191 => 0, 192 => 0, 193 => 0, 194 => 0, 195 => 0, 196 => 0, 197 => 0, 198 => 0, 199 => 1, 200 => 1, 201 => 1, 202 => 1, 203 => 1, 204 => 1, 205 => 1, 206 => 1, 207 => 1, 208 => 1, 209 => 1, 210 => 1, 211 => 1, 212 => 1, 213 => 1, 214 => 1, 215 => 1, 216 => 1, 217 => 1, 218 => 1, 219 => 1, 220 => 1, 221 => 1, 222 
=> 1, 223 => 1, 224 => 1, 225 => 1, 226 => 1, 227 => 1, 228 => 1, 229 => 1, 230 => 1, 231 => 1, 232 => 1, 233 => 1, 234 => 1, 235 => 0, 236 => 0, 237 => 0, 238 => 0, 239 => 0, 240 => 0, 241 => 0, 242 => 0, 243 => 0, 244 => 0, 245 => 0, 246 => 0, 247 => 0, 248 => 0, 249 => 0, 250 => 0, 251 => 0, 252 => 0, 253 => 0, 254 => 0, 255 => 0, 256 => 1, 257 => 1, 258 => 1, 259 => 1, 260 => 1, 261 => 1, 262 => 1, 263 => 1, 264 => 1, 265 => 1, 266 => 1, 267 => 
1, 268 => 1, 269 => 1, 270 => 1, 271 => 1, 272 => 1, 273 => 1, 274 => 1, 275 => 1, 276 => 1, 277 => 1, 278 => 1, 279 => 1, 280 => 1, 281 => 1, 282 => 1, 283 => 1, 284 => 1, 285 => 1, 286 => 1, 287 => 0, 288 => 0, 289 => 0, 290 => 0, 291 => 0, 292 => 0, 293 => 0, 294 => 0, 295 => 0, 296 => 0, 297 => 0, 298 => 0, 299 => 0, 300 => 0, 301 => 1, 302 => 1, 303 => 1, 304 => 1, 305 => 1, 306 => 0, 307 => 0, 308 => 0, 309 => 0, 310 => 0, 311 => 0, 312 => 0, 
313 => 0, 314 => 0, 315 => 0, 316 => 0, 317 => 0, 318 => 0, 319 => 0, 320 => 0, 321 => 0, 322 => 0, 323 => 0, 324 => 0, 325 => 0, 326 => 0, 327 => 0, 328 => 0, 329 => 0, 330 => 0, 331 => 0, 332 => 0, 333 => 1, 334 => 1, 335 => 1, 336 => 1, 337 => 1, 338 => 1, 339 => 1, 340 => 1, 341 => 1, 342 => 1, 343 => 1, 344 => 0, 345 => 0, 346 => 0, 347 => 0, 348 => 0, 349 => 0, 350 => 0, 351 => 0, 352 => 0, 353 => 0, 354 => 0, 355 => 0, 356 => 0, 357 => 0, 358 => 0, 359 => 1, 360 => 1, 361 => 1, 362 => 1, 363 => 1, 364 => 1, 365 => 1, 366 => 1, 367 => 1, 368 => 1, 369 => 1, 370 => 1, 371 => 1, 372 => 1, 373 
=> 1, 374 => 1, 375 => 1, 376 => 1, 377 => 1, 378 => 1, 379 => 1, 380 => 1, 381 => 1, 382 => 1, 383 => 1, 384 => 1, 385 => 1, 386 => 1, 387 => 1, 388 => 1, 389 => 0, 390 => 0, 391 => 0, 392 => 0, 393 => 0, 394 => 0, 395 => 0, 396 => 0, 397 => 1, 398 => 1, 399 => 1, 400 => 1, 401 => 1, 402 => 1, 403 => 1, 404 => 1, 405 => 1, 406 => 1, 407 => 1, 408 => 1, 409 => 1, 410 => 1, 411 => 1, 412 => 1, 413 => 1, 414 => 1, 415 => 1, 416 => 1, 417 => 1, 418 => 
1, 419 => 1, 420 => 1, 421 => 1, 422 => 1, 423 => 1, 424 => 1, 425 => 1, 426 => 1, 427 => 1, 428 => 1, 429 => 1, 430 => 1, 431 => 1, 432 => 1, 433 => 0, 434 => 0, 435 => 0, 436 => 0, 437 => 0, 438 => 0, 439 => 0, 440 => 0, 441 => 0, 442 => 0, 443 => 0, 444 => 0, 445 => 0, 446 => 0, 447 => 0, 448 => 0, 449 => 0, 450 => 0, 451 => 0, 452 => 0, 453 => 0, 454 => 1, 455 => 1, 456 => 1, 457 => 1, 458 => 1, 459 => 1, 460 => 1, 461 => 1, 462 => 1, 463 => 1, 
464 => 1, 465 => 1, 466 => 1, 467 => 1, 468 => 1, 469 => 1, 470 => 1, 471 => 1, 472 => 1, 473 => 1, 474 => 1, 475 => 1, 476 => 1, 477 => 1, 478 => 1, 479 => 1, 480 => 1, 481 => 1, 482 => 1, 483 => 1, 484 => 1, 485 => 0, 486 => 0, 487 => 0, 488 => 0, 489 => 0, 490 => 0, 491 => 0, 492 => 0, 493 => 0, 494 => 0, 495 => 0, 496 => 0, 497 => 0, 498 => 0, 499 => 1, 500 => 1, 501 => 1, 502 => 1, 503 => 1, 504 => 0, 505 => 0, 506 => 0, 507 => 0, 508 => 0, 509 => 0, 510 => 0, 511 => 0, 512 => 0, 513 => 0, 514 => 0, 515 => 0, 516 => 0, 517 => 0, 518 => 0, 519 => 0, 520 => 0, 521 => 0, 522 => 0, 523 => 0, 524 
=> 0, 525 => 0, 526 => 0, 527 => 0, 528 => 0, 529 => 0, 530 => 0, 531 => 1, 532 => 1, 533 => 1, 534 => 1, 535 => 1, 536 => 1, 537 => 1, 538 => 1, 539 => 1, 540 => 1, 541 => 1, 542 => 0, 543 => 0, 544 => 0, 545 => 0, 546 => 0, 547 => 0, 548 => 0, 549 => 0, 550 => 0, 551 => 0, 552 => 0, 553 => 0, 554 => 0, 555 => 0, 556 => 0, 557 => 1, 558 => 1, 559 => 1, 560 => 1, 561 => 1, 562 => 1, 563 => 1, 564 => 1, 565 => 1, 566 => 1, 567 => 1, 568 => 1, 569 => 
1, 570 => 1, 571 => 1, 572 => 1, 573 => 1, 574 => 1, 575 => 1, 576 => 1, 577 => 1, 578 => 1, 579 => 1, 580 => 1, 581 => 1, 582 => 1, 583 => 1, 584 => 1, 585 => 1, 586 => 1, 587 => 0, 588 => 0, 589 => 0, 590 => 0, 591 => 0, 592 => 0, 593 => 0, 594 => 0, 595 => 1, 596 => 1, 597 => 1, 598 => 1, 599 => 1, 600 => 1, 601 => 1, 602 => 1, 603 => 1, 604 => 1, 605 => 1, 606 => 1, 607 => 1, 608 => 1, 609 => 1, 610 => 1, 611 => 1, 612 => 1, 613 => 1, 614 => 1, 
615 => 1, 616 => 1, 617 => 1, 618 => 1, 619 => 1, 620 => 1, 621 => 1, 622 => 1, 623 => 1, 624 => 1, 625 => 1, 626 => 1, 627 => 1, 628 => 1, 629 => 1, 630 => 1, 631 => 0, 632 => 0, 633 => 0, 634 => 0, 635 => 0, 636 => 0, 637 => 0, 638 => 0, 639 => 0, 640 => 0, 641 => 0, 642 => 0, 643 => 0, 644 => 0, 645 => 0, 646 => 0, 647 => 0, 648 => 0, 649 => 0, 650 => 0, 651 => 0, 652 => 1, 653 => 1, 654 => 1, 655 => 1, 656 => 1, 657 => 1, 658 => 1, 659 => 1, 660 => 1, 661 => 1, 662 => 1, 663 => 1, 664 => 1, 665 => 1, 666 => 1, 667 => 1, 668 => 1, 669 => 1, 670 => 1, 671 => 1, 672 => 1, 673 => 1, 674 => 1, 675 
=> 1, 676 => 1, 677 => 1, 678 => 1, 679 => 1, 680 => 1, 681 => 1, 682 => 1, 683 => 0, 684 => 0, 685 => 0, 686 => 0, 687 => 0, 688 => 0, 689 => 0, 690 => 0, 691 => 0, 692 => 0, 693 => 0, 694 => 0, 695 => 0, 696 => 0, 697 => 1, 698 => 1, 699 => 1, 700 => 1, 701 => 1, 702 => 0, 703 => 0, 704 => 0, 705 => 0, 706 => 0, 707 => 0, 708 => 0, 709 => 0, 710 => 0, 711 => 0, 712 => 0, 713 => 0, 714 => 0, 715 => 0, 716 => 0, 717 => 0, 718 => 0, 719 => 0, 720 => 
0, 721 => 0, 722 => 0, 723 => 0, 724 => 0, 725 => 0, 726 => 0, 727 => 0, 728 => 0, 729 => 1, 730 => 1, 731 => 1, 732 => 1, 733 => 1, 734 => 1, 735 => 1, 736 => 1, 737 => 1, 738 => 1, 739 => 1, 740 => 0, 741 => 0, 742 => 0, 743 => 0, 744 => 0, 745 => 0, 746 => 0, 747 => 0, 748 => 0, 749 => 0, 750 => 0, 751 => 0, 752 => 0, 753 => 0, 754 => 0, 755 => 1, 756 => 1, 757 => 1, 758 => 1, 759 => 1, 760 => 1, 761 => 1, 762 => 1, 763 => 1, 764 => 1, 765 => 1, 
766 => 1, 767 => 1, 768 => 1, 769 => 1, 770 => 1, 771 => 1, 772 => 1, 773 => 1, 774 => 1, 775 => 1, 776 => 1, 777 => 1, 778 => 1, 779 => 1, 780 => 1, 781 => 1, 782 => 1, 783 => 1, 784 => 1, 785 => 0, 786 => 0, 787 => 0, 788 => 0, 789 => 0, 790 => 0, 791 => 0, 792 => 0, 793 => 1, 794 => 1, 795 => 1, 796 => 1, 797 => 1, 798 => 1, 799 => 1, 800 => 1, 801 => 1, 802 => 1, 803 => 1, 804 => 1, 805 => 1, 806 => 1, 807 => 1, 808 => 1, 809 => 1, 810 => 1, 811 => 1, 812 => 1, 813 => 1, 814 => 1, 815 => 1, 816 => 1, 817 => 1, 818 => 1, 819 => 1, 820 => 1, 821 => 1, 822 => 1, 823 => 1, 824 => 1, 825 => 1, 826 
=> 1, 827 => 1, 828 => 1, 829 => 0, 830 => 0, 831 => 0, 832 => 0, 833 => 0, 834 => 0, 835 => 0, 836 => 0, 837 => 0, 838 => 0, 839 => 0, 840 => 0, 841 => 0, 842 => 0, 843 => 0, 844 => 0, 845 => 0, 846 => 0, 847 => 0, 848 => 0, 849 => 0, 850 => 1, 851 => 1, 852 => 1, 853 => 1, 854 => 1, 855 => 1, 856 => 1, 857 => 1, 858 => 1, 859 => 1, 860 => 1, 861 => 1, 862 => 1, 863 => 1, 864 => 1, 865 => 1, 866 => 1, 867 => 1, 868 => 1, 869 => 1, 870 => 1, 871 => 
1, 872 => 1, 873 => 1, 874 => 1, 875 => 1, 876 => 1, 877 => 1, 878 => 1, 879 => 1, 880 => 1, 881 => 0, 882 => 0, 883 => 0, 884 => 0, 885 => 0, 886 => 0, 887 => 0, 888 => 0, 889 => 0, 890 => 0, 891 => 0, 892 => 0, 893 => 0, 894 => 0, 895 => 1, 896 => 1, 897 => 1, 898 => 1, 899 => 1, 900 => 0, 901 => 0, 902 => 0, 903 => 0, 904 => 0, 905 => 0, 906 => 0, 907 => 0, 908 => 0, 909 => 0, 910 => 0, 911 => 0, 912 => 0, 913 => 0, 914 => 0, 915 => 0, 916 => 0, 
917 => 0, 918 => 0, 919 => 0, 920 => 0, 921 => 0, 922 => 0, 923 => 0, 924 => 0, 925 => 0, 926 => 0, 927 => 1, 928 => 1, 929 => 1, 930 => 1, 931 => 1, 932 => 1, 933 => 1, 934 => 1, 935 => 1, 936 => 1, 937 => 1, 938 => 0, 939 => 0, 940 => 0, 941 => 0, 942 => 0, 943 => 0, 944 => 0, 945 => 0, 946 => 0, 947 => 0, 948 => 0, 949 => 0, 950 => 0, 951 => 0, 952 => 0, 953 => 1, 954 => 1, 955 => 1, 956 => 1, 957 => 1, 958 => 1, 959 => 1, 960 => 1, 961 => 1, 962 => 1, 963 => 1, 964 => 1, 965 => 1, 966 => 1, 967 => 1, 968 => 1, 969 => 1, 970 => 1, 971 => 1, 972 => 1, 973 => 1, 974 => 1, 975 => 1, 976 => 1, 977 
=> 1, 978 => 1, 979 => 1, 980 => 1, 981 => 1, 982 => 1, 983 => 0, 984 => 0, 985 => 0, 986 => 0, 987 => 0, 988 => 0, 989 => 0, 990 => 0, 991 => 1, 992 => 1, 993 => 1, 994 => 1, 995 => 1, 996 => 1, 997 => 1, 998 => 1, 999 => 1, 1000 => 1, 1001 => 1, 1002 => 1, 1003 => 1, 1004 => 1, 1005 => 1, 1006 => 1, 1007 => 1, 1008 => 1, 1009 => 1, 1010 => 1, 1011 => 1, 1012 => 1, 1013 => 1, 1014 => 1, 1015 => 1, 1016 => 1, 1017 => 1, 1018 => 1, 1019 => 1, 1020 => 1, 1021 => 1, 1022 => 1, 1023 => 1, 1024 => 1, 1025 => 1, 1026 => 1, 1027 => 0, 1028 => 0, 1029 => 0, 1030 => 0, 1031 => 0, 1032 => 0, 1033 => 0, 1034 => 0, 1035 => 0, 1036 => 0, 1037 => 0, 1038 => 0, 1039 => 0, 1040 => 0, 1041 => 0, 1042 => 0, 1043 => 0, 1044 => 0, 1045 => 0, 1046 => 0, 1047 => 0, 1048 => 1, 1049 => 1, 1050 => 1, 1051 => 1, 1052 => 1, 1053 => 1, 1054 => 1, 1055 => 1, 1056 => 1, 1057 => 1, 1058 => 1, 1059 => 1, 1060 => 1, 1061 => 1, 1062 => 1, 1063 => 1, 1064 => 1, 1065 => 1, 1066 => 1, 1067 => 1, 1068 => 1, 1069 => 1, 1070 => 1, 1071 => 1, 1072 => 1, 1073 => 1, 1074 => 1, 1075 => 1, 1076 => 1, 1077 => 1, 1078 => 1, 1079 => 0, 1080 => 0, 1081 => 0, 1082 => 0, 1083 => 0, 1084 => 0, 1085 => 0, 1086 => 0, 1087 => 0, 1088 => 0, 1089 => 0, 1090 => 0, 1091 => 0, 1092 => 0, 1093 => 1, 1094 => 1, 1095 => 1, 1096 => 1, 1097 => 1, 1098 => 0, 1099 => 0, 1100 => 0, 1101 => 0, 1102 => 0, 
1103 => 0, 1104 => 0, 1105 => 0, 1106 => 0, 1107 => 0, 1108 => 0, 1109 => 0, 1110 => 0, 1111 => 0, 1112 => 0, 1113 => 0, 1114 => 0, 1115 => 0, 1116 => 
0, 1117 => 0, 1118 => 0, 1119 => 0, 1120 => 0, 1121 => 0, 1122 => 0, 1123 => 0, 1124 => 0, 1125 => 1, 1126 => 1, 1127 => 1, 1128 => 1, 1129 => 1, 1130 
=> 1, 1131 => 1, 1132 => 1, 1133 => 1, 1134 => 1, 1135 => 1, 1136 => 0, 1137 => 0, 1138 => 0, 1139 => 0, 1140 => 0, 1141 => 0, 1142 => 0, 1143 => 0, 1144 => 0, 1145 => 0, 1146 => 0, 1147 => 0, 1148 => 0, 1149 => 0, 1150 => 0, 1151 => 1, 1152 => 1, 1153 => 1, 1154 => 1, 1155 => 1, 1156 => 1, 1157 => 1, 1158 => 1, 1159 => 1, 1160 => 1, 1161 => 1, 1162 => 1, 1163 => 1, 1164 => 1, 1165 => 1, 1166 => 1, 1167 => 1, 1168 => 1, 1169 => 1, 1170 => 1, 1171 => 1, 1172 => 1, 1173 => 1, 1174 => 1, 1175 => 1, 1176 => 1, 1177 => 1, 1178 => 1, 1179 => 1, 1180 => 1, 1181 => 0, 1182 => 0, 1183 => 0, 1184 => 0, 1185 => 0, 1186 => 0, 1187 => 0, 1188 => 0, 1189 => 1, 1190 => 1, 1191 => 1, 1192 => 1, 1193 => 1, 1194 => 1, 1195 => 1, 1196 => 1, 1197 => 1, 1198 => 1, 1199 => 1, 1200 => 0, 1201 => 0, 1202 => 0, 1203 => 0, 1204 => 0, 1205 => 0, 1206 => 0, 1207 => 0, 1208 => 0, 1209 => 0, 1210 => 0, 1211 => 0, 1212 => 0, 1213 => 0, 1214 => 0, 1215 => 0, 1216 => 0, 1217 => 0, 1218 => 0, 1219 => 0, 1220 => 0, 1221 => 1, 1222 => 1, 1223 => 1, 1224 => 1, 1225 => 1, 1226 => 0, 1227 => 0, 1228 => 0, 1229 => 0, 1230 => 0, 1231 => 0, 1232 => 0, 1233 => 0, 1234 => 0, 1235 => 0, 1236 => 0, 1237 => 0, 1238 => 0, 1239 => 0, 1240 => 0, 1241 => 0, 1242 => 0, 1243 => 0, 1244 => 0, 1245 => 0, 1246 => 1, 1247 => 1, 1248 => 1, 1249 => 1, 1250 => 1, 1251 => 0, 1252 => 0, 1253 => 0, 
1254 => 0, 1255 => 0, 1256 => 0, 1257 => 0, 1258 => 0, 1259 => 0, 1260 => 0, 1261 => 0, 1262 => 0, 1263 => 0, 1264 => 0, 1265 => 0, 1266 => 0, 1267 => 
0, 1268 => 0, 1269 => 0, 1270 => 0, 1271 => 0, 1272 => 1, 1273 => 1, 1274 => 1, 1275 => 1, 1276 => 1, 1277 => 0, 1278 => 0, 1279 => 0, 1280 => 0, 1281 
=> 0, 1282 => 0, 1283 => 0, 1284 => 0, 1285 => 0, 1286 => 0, 1287 => 0, 1288 => 0, 1289 => 0, 1290 => 0, 1291 => 1, 1292 => 1, 1293 => 1, 1294 => 1, 1295 => 1, 1296 => 0, 1297 => 0, 1298 => 0, 1299 => 0, 1300 => 0, 1301 => 0, 1302 => 0, 1303 => 0, 1304 => 0, 1305 => 0, 1306 => 0, 1307 => 0, 1308 => 0, 1309 => 0, 1310 => 0, 1311 => 0, 1312 => 0, 1313 => 0, 1314 => 0, 1315 => 0, 1316 => 0, 1317 => 0, 1318 => 0, 1319 => 0, 1320 => 0, 1321 => 0, 1322 => 0, 1323 => 1, 1324 => 1, 1325 => 1, 1326 => 1, 1327 => 1, 1328 => 1, 1329 => 1, 1330 => 1, 1331 => 1, 1332 => 1, 1333 => 1, 1334 => 0, 1335 => 0, 1336 => 0, 1337 => 0, 1338 => 0, 1339 => 0, 1340 => 0, 1341 => 0, 1342 => 0, 1343 => 0, 1344 => 0, 1345 => 0, 1346 => 0, 1347 => 0, 1348 => 1, 1349 => 1, 1350 => 1, 1351 => 1, 1352 => 1, 1353 => 0, 1354 => 0, 1355 => 0, 1356 => 0, 1357 => 0, 1358 => 0, 1359 => 0, 1360 => 0, 1361 => 0, 1362 => 0, 1363 => 0, 1364 => 0, 1365 => 0, 1366 => 0, 1367 => 0, 1368 => 0, 1369 => 0, 1370 => 0, 1371 => 0, 1372 => 0, 1373 => 0, 1374 => 1, 1375 => 1, 1376 => 1, 1377 => 1, 1378 => 1, 1379 => 0, 1380 => 0, 1381 => 0, 1382 => 0, 1383 => 0, 1384 => 0, 1385 => 0, 1386 => 0, 1387 => 1, 1388 => 1, 1389 => 1, 1390 => 1, 1391 => 1, 1392 => 1, 1393 => 1, 1394 => 1, 1395 => 1, 1396 => 1, 1397 => 1, 1398 => 0, 1399 => 0, 1400 => 0, 1401 => 0, 1402 => 0, 1403 => 0, 1404 => 0, 
1405 => 0, 1406 => 0, 1407 => 0, 1408 => 0, 1409 => 0, 1410 => 0, 1411 => 0, 1412 => 0, 1413 => 0, 1414 => 0, 1415 => 0, 1416 => 0, 1417 => 0, 1418 => 
0, 1419 => 1, 1420 => 1, 1421 => 1, 1422 => 1, 1423 => 1, 1424 => 1, 1425 => 1, 1426 => 1, 1427 => 1, 1428 => 1, 1429 => 1, 1430 => 0, 1431 => 0, 1432 
=> 0, 1433 => 0, 1434 => 0, 1435 => 0, 1436 => 0, 1437 => 0, 1438 => 1, 1439 => 1, 1440 => 1, 1441 => 1, 1442 => 1, 1443 => 1, 1444 => 1, 1445 => 1, 1446 => 1, 1447 => 1, 1448 => 1, 1449 => 0, 1450 => 0, 1451 => 0, 1452 => 0, 1453 => 0, 1454 => 0, 1455 => 0, 1456 => 0, 1457 => 0, 1458 => 0, 1459 => 0, 1460 => 0, 1461 => 0, 1462 => 0, 1463 => 0, 1464 => 0, 1465 => 0, 1466 => 0, 1467 => 0, 1468 => 0, 1469 => 0, 1470 => 1, 1471 => 1, 1472 => 1, 1473 => 1, 1474 => 1, 1475 => 1, 1476 => 1, 1477 => 1, 1478 => 1, 1479 => 1, 1480 => 1, 1481 => 0, 1482 => 0, 1483 => 0, 1484 => 0, 1485 => 0, 1486 => 0, 1487 => 0, 1488 => 0, 1489 => 1, 1490 => 1, 1491 => 1, 1492 => 1, 1493 => 1, 1494 => 1, 1495 => 1, 1496 => 1, 1497 => 1, 1498 => 1, 1499 => 1, 1500 => 0, 1501 => 0, 1502 => 0, 1503 => 0, 1504 => 0, 1505 => 0, 1506 => 0, 1507 => 0, 1508 => 0, 1509 => 0, 1510 => 0, 1511 => 0, 1512 => 0, 1513 => 0, 1514 => 0, 1515 => 0, 1516 => 0, 1517 => 0, 1518 => 0, 1519 => 0, 1520 => 0, 1521 => 1, 1522 => 1, 1523 => 1, 1524 => 1, 1525 => 1, 1526 => 1, 1527 => 1, 1528 => 1, 1529 => 1, 1530 => 1, 1531 => 1, 1532 => 0, 1533 => 0, 1534 => 0, 1535 => 0, 1536 => 0, 1537 => 0, 1538 => 0, 1539 => 0, 1540 => 1, 1541 => 1, 1542 => 1, 1543 => 1, 1544 => 1, 1545 => 1, 1546 => 1, 1547 => 1, 1548 => 1, 1549 => 1, 1550 => 1, 1551 => 0, 1552 => 0, 1553 => 0, 1554 => 0, 1555 => 0, 
1556 => 0, 1557 => 0, 1558 => 0, 1559 => 0, 1560 => 0, 1561 => 0, 1562 => 0, 1563 => 0, 1564 => 0, 1565 => 0, 1566 => 0, 1567 => 0, 1568 => 0, 1569 => 
0, 1570 => 0, 1571 => 0, 1572 => 1, 1573 => 1, 1574 => 1, 1575 => 1, 1576 => 1, 1577 => 1, 1578 => 1, 1579 => 1, 1580 => 1, 1581 => 1, 1582 => 1, 1583 
=> 0, 1584 => 0, 1585 => 1, 1586 => 1, 1587 => 1, 1588 => 1, 1589 => 1, 1590 => 1, 1591 => 1, 1592 => 1, 1593 => 1, 1594 => 1, 1595 => 1, 1596 => 0, 1597 => 0, 1598 => 0, 1599 => 0, 1600 => 0, 1601 => 0, 1602 => 0, 1603 => 0, 1604 => 0, 1605 => 0, 1606 => 0, 1607 => 0, 1608 => 0, 1609 => 0, 1610 => 0, 1611 => 0, 1612 => 0, 1613 => 0, 1614 => 0, 1615 => 0, 1616 => 0, 1617 => 1, 1618 => 1, 1619 => 1, 1620 => 1, 1621 => 1, 1622 => 1, 1623 => 1, 1624 => 1, 1625 => 1, 1626 => 1, 1627 => 1, 1628 => 0, 1629 => 0, 1630 => 0, 1631 => 0, 1632 => 0, 1633 => 0, 1634 => 0, 1635 => 0, 1636 => 1, 1637 => 1, 1638 => 1, 1639 => 1, 1640 => 1, 1641 => 1, 1642 => 1, 1643 => 1, 1644 => 1, 1645 => 1, 1646 => 1, 1647 => 0, 1648 => 0, 1649 => 0, 1650 => 0, 1651 => 0, 1652 => 0, 1653 => 0, 1654 => 0, 1655 => 0, 1656 => 0, 1657 => 0, 1658 => 0, 1659 => 0, 1660 => 0, 1661 => 0, 1662 => 0, 1663 => 0, 1664 => 0, 1665 => 0, 1666 => 0, 1667 => 0, 1668 => 1, 1669 => 1, 1670 => 1, 1671 => 1, 1672 => 1, 1673 => 1, 1674 => 1, 1675 => 1, 1676 => 1, 1677 => 1, 1678 => 1, 1679 => 0, 1680 => 0, 1681 => 0, 1682 => 0, 1683 => 0, 1684 => 0, 1685 => 0, 1686 => 0, 1687 => 1, 1688 => 1, 1689 => 1, 1690 => 1, 1691 => 1, 1692 => 1, 1693 => 1, 1694 => 1, 1695 => 1, 1696 => 1, 1697 => 1, 1698 => 0, 1699 => 0, 1700 => 0, 1701 => 0, 1702 => 0, 1703 => 0, 1704 => 0, 1705 => 0, 1706 => 0, 
1707 => 0, 1708 => 0, 1709 => 0, 1710 => 0, 1711 => 0, 1712 => 0, 1713 => 0, 1714 => 0, 1715 => 0, 1716 => 0, 1717 => 0, 1718 => 0, 1719 => 1, 1720 => 
1, 1721 => 1, 1722 => 1, 1723 => 1, 1724 => 1, 1725 => 1, 1726 => 1, 1727 => 1, 1728 => 1, 1729 => 1, 1730 => 0, 1731 => 0, 1732 => 0, 1733 => 0, 1734 
=> 0, 1735 => 0, 1736 => 0, 1737 => 0, 1738 => 1, 1739 => 1, 1740 => 1, 1741 => 1, 1742 => 1, 1743 => 1, 1744 => 1, 1745 => 1, 1746 => 1, 1747 => 1, 1748 => 1, 1749 => 0, 1750 => 0, 1751 => 0, 1752 => 0, 1753 => 0, 1754 => 0, 1755 => 0, 1756 => 0, 1757 => 0, 1758 => 0, 1759 => 0, 1760 => 0, 1761 => 0, 1762 => 0, 1763 => 0, 1764 => 0, 1765 => 0, 1766 => 0, 1767 => 0, 1768 => 0, 1769 => 0, 1770 => 1, 1771 => 1, 1772 => 1, 1773 => 1, 1774 => 1, 1775 => 1, 1776 => 1, 1777 => 1, 1778 => 1, 1779 => 1, 1780 => 1, 1781 => 0, 1782 => 0, 1783 => 1, 1784 => 1, 1785 => 1, 1786 => 1, 1787 => 1, 1788 => 1, 1789 => 1, 1790 => 1, 1791 => 1, 1792 => 1, 1793 => 1, 1794 => 0, 1795 => 0, 1796 => 0, 1797 => 0, 1798 => 0, 1799 => 0, 1800 => 0, 1801 => 0, 1802 => 0, 1803 => 0, 1804 => 0, 1805 => 0, 1806 => 0, 1807 => 0, 1808 => 0, 1809 => 0, 1810 => 0, 1811 => 0, 1812 => 0, 1813 => 0, 1814 => 0, 1815 => 1, 1816 => 1, 1817 => 1, 1818 => 1, 1819 => 1, 1820 => 1, 1821 => 1, 1822 => 1, 1823 => 1, 1824 => 1, 1825 => 1, 1826 => 0, 1827 => 0, 1828 => 0, 1829 => 0, 1830 => 0, 1831 => 0, 1832 => 0, 1833 => 0, 1834 => 1, 1835 => 1, 1836 => 1, 1837 => 1, 1838 => 1, 1839 => 1, 1840 => 1, 1841 => 1, 1842 => 1, 1843 => 1, 1844 => 1, 1845 => 0, 1846 => 0, 1847 => 0, 1848 => 0, 1849 => 0, 1850 => 0, 1851 => 0, 1852 => 0, 1853 => 0, 1854 => 0, 1855 => 0, 1856 => 0, 1857 => 0, 
1858 => 0, 1859 => 0, 1860 => 0, 1861 => 0, 1862 => 0, 1863 => 0, 1864 => 0, 1865 => 0, 1866 => 1, 1867 => 1, 1868 => 1, 1869 => 1, 1870 => 1, 1871 => 
1, 1872 => 1, 1873 => 1, 1874 => 1, 1875 => 1, 1876 => 1, 1877 => 0, 1878 => 0, 1879 => 0, 1880 => 0, 1881 => 0, 1882 => 0, 1883 => 0, 1884 => 0, 1885 
=> 1, 1886 => 1, 1887 => 1, 1888 => 1, 1889 => 1, 1890 => 1, 1891 => 1, 1892 => 1, 1893 => 1, 1894 => 1, 1895 => 1, 1896 => 0, 1897 => 0, 1898 => 0, 1899 => 0, 1900 => 0, 1901 => 0, 1902 => 0, 1903 => 0, 1904 => 0, 1905 => 0, 1906 => 0, 1907 => 0, 1908 => 0, 1909 => 0, 1910 => 0, 1911 => 0, 1912 => 0, 1913 => 0, 1914 => 0, 1915 => 0, 1916 => 0, 1917 => 1, 1918 => 1, 1919 => 1, 1920 => 1, 1921 => 1, 1922 => 1, 1923 => 1, 1924 => 1, 1925 => 1, 1926 => 1, 1927 => 1, 1928 => 0, 1929 => 0, 1930 => 0, 1931 => 0, 1932 => 0, 1933 => 0, 1934 => 0, 1935 => 0, 1936 => 1, 1937 => 1, 1938 => 1, 1939 => 1, 1940 => 1, 1941 => 1, 1942 => 1, 1943 => 1, 1944 => 1, 1945 => 1, 1946 => 1, 1947 => 0, 1948 => 0, 1949 => 0, 1950 => 0, 1951 => 0, 1952 => 0, 1953 => 0, 1954 => 0, 1955 => 0, 1956 => 0, 1957 => 0, 1958 => 0, 1959 => 0, 1960 => 0, 1961 => 0, 1962 => 0, 1963 => 0, 1964 => 0, 1965 => 0, 1966 => 0, 1967 => 0, 1968 => 1, 1969 => 1, 1970 => 1, 1971 => 1, 1972 => 1, 1973 => 1, 1974 => 1, 1975 => 1, 1976 => 1, 1977 => 1, 1978 => 1, 1979 => 0, 1980 => 0, 1981 => 1, 1982 => 1, 1983 => 1, 1984 => 1, 1985 => 1, 1986 => 1, 1987 => 1, 1988 => 1, 1989 => 1, 1990 => 1, 1991 => 1, 1992 => 0, 1993 => 0, 1994 => 0, 1995 => 0, 1996 => 0, 1997 => 0, 1998 => 0, 1999 => 0, 2000 => 0, 2001 => 0, 2002 => 0, 2003 => 0, 2004 => 0, 2005 => 0, 2006 => 0, 2007 => 0, 2008 => 0, 
2009 => 0, 2010 => 0, 2011 => 0, 2012 => 0, 2013 => 1, 2014 => 1, 2015 => 1, 2016 => 1, 2017 => 1, 2018 => 1, 2019 => 1, 2020 => 1, 2021 => 1, 2022 => 
1, 2023 => 1, 2024 => 0, 2025 => 0, 2026 => 0, 2027 => 0, 2028 => 0, 2029 => 0, 2030 => 0, 2031 => 0, 2032 => 1, 2033 => 1, 2034 => 1, 2035 => 1, 2036 
=> 1, 2037 => 1, 2038 => 1, 2039 => 1, 2040 => 1, 2041 => 1, 2042 => 1, 2043 => 0, 2044 => 0, 2045 => 0, 2046 => 0, 2047 => 0, 2048 => 0, 2049 => 0, 2050 => 0, 2051 => 0, 2052 => 0, 2053 => 0, 2054 => 0, 2055 => 0, 2056 => 0, 2057 => 0, 2058 => 0, 2059 => 0, 2060 => 0, 2061 => 0, 2062 => 0, 2063 => 0, 2064 => 1, 2065 => 1, 2066 => 1, 2067 => 1, 2068 => 1, 2069 => 1, 2070 => 1, 2071 => 1, 2072 => 1, 2073 => 1, 2074 => 1, 2075 => 0, 2076 => 0, 2077 => 0, 2078 => 0, 2079 => 0, 2080 => 0, 2081 => 0, 2082 => 0, 2083 => 1, 2084 => 1, 2085 => 1, 2086 => 1, 2087 => 1, 2088 => 1, 2089 => 1, 2090 => 1, 2091 => 1, 2092 => 1, 2093 => 1, 2094 => 0, 2095 => 0, 2096 => 0, 2097 => 0, 2098 => 0, 2099 => 0, 2100 => 0, 2101 => 0, 2102 => 0, 2103 => 0, 2104 => 0, 2105 => 0, 2106 => 0, 2107 => 0, 2108 => 0, 2109 => 0, 2110 => 0, 2111 => 0, 2112 => 0, 2113 => 0, 2114 => 0, 2115 => 1, 2116 => 1, 2117 => 1, 2118 => 1, 2119 => 1, 2120 => 1, 2121 => 1, 2122 => 1, 2123 => 1, 2124 => 1, 2125 => 1, 2126 => 0, 2127 => 0, 2128 => 0, 2129 => 0, 2130 => 0, 2131 => 0, 2132 => 0, 2133 => 0, 2134 => 1, 2135 => 1, 2136 => 1, 2137 => 1, 2138 => 1, 2139 => 1, 2140 => 1, 2141 => 1, 2142 => 1, 2143 => 1, 2144 => 1, 2145 => 0, 2146 => 0, 2147 => 0, 2148 => 0, 2149 => 0, 2150 => 0, 2151 => 0, 2152 => 0, 2153 => 0, 2154 => 0, 2155 => 0, 2156 => 0, 2157 => 0, 2158 => 0, 2159 => 0, 
2160 => 0, 2161 => 0, 2162 => 0, 2163 => 0, 2164 => 0, 2165 => 0, 2166 => 1, 2167 => 1, 2168 => 1, 2169 => 1, 2170 => 1, 2171 => 1, 2172 => 1, 2173 => 
1, 2174 => 1, 2175 => 1, 2176 => 1, 2177 => 0, 2178 => 0, 2179 => 1, 2180 => 1, 2181 => 1, 2182 => 1, 2183 => 1, 2184 => 1, 2185 => 1, 2186 => 1, 2187 
=> 1, 2188 => 1, 2189 => 1, 2190 => 0, 2191 => 0, 2192 => 0, 2193 => 0, 2194 => 0, 2195 => 0, 2196 => 0, 2197 => 0, 2198 => 0, 2199 => 0, 2200 => 0, 2201 => 0, 2202 => 0, 2203 => 0, 2204 => 0, 2205 => 0, 2206 => 0, 2207 => 0, 2208 => 0, 2209 => 0, 2210 => 0, 2211 => 1, 2212 => 1, 2213 => 1, 2214 => 1, 2215 => 1, 2216 => 1, 2217 => 1, 2218 => 1, 2219 => 1, 2220 => 1, 2221 => 1, 2222 => 0, 2223 => 0, 2224 => 0, 2225 => 0, 2226 => 0, 2227 => 0, 2228 => 0, 2229 => 0, 2230 => 1, 2231 => 1, 2232 => 1, 2233 => 1, 2234 => 1, 2235 => 1, 2236 => 1, 2237 => 1, 2238 => 1, 2239 => 1, 2240 => 1, 2241 => 0, 2242 => 0, 2243 => 0, 2244 => 0, 2245 => 0, 2246 => 0, 2247 => 0, 2248 => 0, 2249 => 0, 2250 => 0, 2251 => 0, 2252 => 0, 2253 => 0, 2254 => 0, 2255 => 0, 2256 => 0, 2257 => 0, 2258 => 0, 2259 => 0, 2260 => 0, 2261 => 0, 2262 => 1, 2263 => 1, 2264 => 1, 2265 => 1, 2266 => 1, 2267 => 1, 2268 => 1, 2269 => 1, 2270 => 1, 2271 => 1, 2272 => 1, 2273 => 0, 2274 => 0, 2275 => 0, 2276 => 0, 2277 => 0, 2278 => 0, 2279 => 0, 2280 => 0, 2281 => 1, 2282 => 1, 2283 => 1, 2284 => 1, 2285 => 1, 2286 => 1, 2287 => 1, 2288 => 1, 2289 => 1, 2290 => 1, 2291 => 1, 2292 => 0, 2293 => 0, 2294 => 0, 2295 => 0, 2296 => 0, 2297 => 0, 2298 => 0, 2299 => 0, 2300 => 0, 2301 => 0, 2302 => 0, 2303 => 0, 2304 => 0, 2305 => 0, 2306 => 0, 2307 => 0, 2308 => 0, 2309 => 0, 2310 => 0, 
2311 => 0, 2312 => 0, 2313 => 1, 2314 => 1, 2315 => 1, 2316 => 1, 2317 => 1, 2318 => 1, 2319 => 1, 2320 => 1, 2321 => 1, 2322 => 1, 2323 => 1, 2324 => 
0, 2325 => 0, 2326 => 0, 2327 => 0, 2328 => 0, 2329 => 0, 2330 => 0, 2331 => 0, 2332 => 1, 2333 => 1, 2334 => 1, 2335 => 1, 2336 => 1, 2337 => 1, 2338 
=> 1, 2339 => 1, 2340 => 1, 2341 => 1, 2342 => 1, 2343 => 0, 2344 => 0, 2345 => 0, 2346 => 0, 2347 => 0, 2348 => 0, 2349 => 0, 2350 => 0, 2351 => 0, 2352 => 0, 2353 => 0, 2354 => 0, 2355 => 0, 2356 => 0, 2357 => 0, 2358 => 0, 2359 => 0, 2360 => 0, 2361 => 0, 2362 => 0, 2363 => 0, 2364 => 1, 2365 => 1, 2366 => 1, 2367 => 1, 2368 => 1, 2369 => 1, 2370 => 1, 2371 => 1, 2372 => 1, 2373 => 1, 2374 => 1, 2375 => 0, 2376 => 0, 2377 => 1, 2378 => 1, 2379 => 1, 2380 => 1, 2381 => 1, 2382 => 1, 2383 => 1, 2384 => 1, 2385 => 1, 2386 => 1, 2387 => 1, 2388 => 0, 2389 => 0, 2390 => 0, 2391 => 0, 2392 => 0, 2393 => 0, 2394 => 0, 2395 => 0, 2396 => 0, 2397 => 0, 2398 => 0, 2399 => 0, 2400 => 0, 2401 => 0, 2402 => 0, 2403 => 0, 2404 => 0, 2405 => 0, 2406 => 0, 2407 => 0, 2408 => 0, 2409 => 1, 2410 => 1, 2411 => 1, 2412 => 1, 2413 => 1, 2414 => 1, 2415 => 1, 2416 => 1, 2417 => 1, 2418 => 1, 2419 => 1, 2420 => 0, 2421 => 0, 2422 => 0, 2423 => 0, 2424 => 0, 2425 => 0, 2426 => 0, 2427 => 0, 2428 => 1, 2429 => 1, 2430 => 1, 2431 => 1, 2432 => 1, 2433 => 1, 2434 => 1, 2435 => 1, 2436 => 1, 2437 => 1, 2438 => 1, 2439 => 0, 2440 => 0, 2441 => 0, 2442 => 0, 2443 => 0, 2444 => 0, 2445 => 0, 2446 => 0, 2447 => 0, 2448 => 0, 2449 => 0, 2450 => 0, 2451 => 0, 2452 => 0, 2453 => 0, 2454 => 0, 2455 => 0, 2456 => 0, 2457 => 0, 2458 => 0, 2459 => 0, 2460 => 1, 2461 => 1, 
2462 => 1, 2463 => 1, 2464 => 1, 2465 => 1, 2466 => 1, 2467 => 1, 2468 => 1, 2469 => 1, 2470 => 1, 2471 => 0, 2472 => 0, 2473 => 0, 2474 => 0, 2475 => 
0, 2476 => 0, 2477 => 0, 2478 => 0, 2479 => 1, 2480 => 1, 2481 => 1, 2482 => 1, 2483 => 1, 2484 => 1, 2485 => 1, 2486 => 1, 2487 => 1, 2488 => 1, 2489 
=> 1, 2490 => 0, 2491 => 0, 2492 => 0, 2493 => 0, 2494 => 0, 2495 => 0, 2496 => 0, 2497 => 0, 2498 => 0, 2499 => 0, 2500 => 0, 2501 => 0, 2502 => 0, 2503 => 0, 2504 => 0, 2505 => 0, 2506 => 0, 2507 => 0, 2508 => 0, 2509 => 0, 2510 => 0, 2511 => 1, 2512 => 1, 2513 => 1, 2514 => 1, 2515 => 1, 2516 => 1, 2517 => 1, 2518 => 1, 2519 => 1, 2520 => 1, 2521 => 1, 2522 => 0, 2523 => 0, 2524 => 0, 2525 => 0, 2526 => 0, 2527 => 0, 2528 => 0, 2529 => 0, 2530 => 1, 2531 => 1, 2532 => 1, 2533 => 1, 2534 => 1, 2535 => 1, 2536 => 1, 2537 => 1, 2538 => 1, 2539 => 1, 2540 => 1, 2541 => 0, 2542 => 0, 2543 => 0, 2544 => 0, 2545 => 0, 2546 => 0, 2547 => 0, 2548 => 0, 2549 => 0, 2550 => 0, 2551 => 0, 2552 => 0, 2553 => 0, 2554 => 0, 2555 => 0, 2556 => 0, 2557 => 0, 2558 => 0, 2559 => 0, 2560 => 0, 2561 => 0, 2562 => 0, 2563 => 0, 2564 => 0, 2565 => 0, 2566 => 0, 2567 => 0, 2568 => 0, 2569 => 0, 2570 => 0, 2571 => 0, 2572 => 0, 2573 => 0, 2574 => 0, 2575 => 1, 2576 => 1, 2577 => 1, 2578 => 1, 2579 => 1, 2580 => 1, 2581 => 1, 2582 => 1, 2583 => 1, 2584 => 1, 2585 => 1, 2586 => 0, 2587 => 0, 2588 => 0, 2589 => 0, 2590 => 0, 2591 => 0, 2592 => 0, 2593 => 0, 2594 => 0, 2595 => 0, 2596 => 0, 2597 => 0, 2598 => 0, 2599 => 0, 2600 => 0, 2601 => 0, 2602 => 0, 2603 => 0, 2604 => 0, 2605 => 0, 2606 => 0, 2607 => 1, 2608 => 1, 2609 => 1, 2610 => 1, 2611 => 1, 2612 => 1, 
2613 => 1, 2614 => 1, 2615 => 1, 2616 => 1, 2617 => 1, 2618 => 0, 2619 => 0, 2620 => 0, 2621 => 0, 2622 => 0, 2623 => 0, 2624 => 0, 2625 => 0, 2626 => 
1, 2627 => 1, 2628 => 1, 2629 => 1, 2630 => 1, 2631 => 1, 2632 => 1, 2633 => 1, 2634 => 1, 2635 => 1, 2636 => 1, 2637 => 0, 2638 => 0, 2639 => 0, 2640 
=> 0, 2641 => 0, 2642 => 0, 2643 => 0, 2644 => 0, 2645 => 0, 2646 => 0, 2647 => 0, 2648 => 0, 2649 => 0, 2650 => 0, 2651 => 0, 2652 => 0, 2653 => 0, 2654 => 0, 2655 => 0, 2656 => 0, 2657 => 0, 2658 => 1, 2659 => 1, 2660 => 1, 2661 => 1, 2662 => 1, 2663 => 1, 2664 => 1, 2665 => 1, 2666 => 1, 2667 => 1, 2668 => 1, 2669 => 0, 2670 => 0, 2671 => 0, 2672 => 0, 2673 => 0, 2674 => 0, 2675 => 0, 2676 => 0, 2677 => 1, 2678 => 1, 2679 => 1, 2680 => 1, 2681 => 1, 2682 => 1, 2683 => 1, 2684 => 1, 2685 => 1, 2686 => 1, 2687 => 1, 2688 => 1, 2689 => 0, 2690 => 0, 2691 => 0, 2692 => 0, 2693 => 0, 2694 => 1, 2695 => 0, 2696 => 0, 2697 => 0, 2698 => 0, 2699 => 0, 2700 => 0, 2701 => 0, 2702 => 0, 2703 => 0, 2704 => 0, 2705 => 0, 2706 => 0, 2707 => 0, 2708 => 0, 2709 => 1, 2710 => 1, 2711 => 1, 2712 => 1, 2713 => 1, 2714 => 1, 2715 => 1, 2716 => 1, 2717 => 1, 2718 => 1, 2719 => 1, 2720 => 0, 2721 => 0, 2722 => 0, 2723 => 0, 2724 => 0, 2725 => 0, 2726 => 0, 2727 => 0, 2728 => 1, 2729 => 1, 2730 => 1, 2731 => 1, 2732 => 1, 2733 => 1, 2734 => 1, 2735 => 1, 2736 => 1, 2737 => 1, 2738 => 1, 2739 => 0, 2740 => 0, 2741 => 0, 2742 => 0, 2743 => 0, 2744 => 0, 2745 => 0, 2746 => 0, 2747 => 0, 2748 => 0, 2749 => 0, 2750 => 0, 2751 => 0, 2752 => 0, 2753 => 0, 2754 => 0, 2755 => 0, 2756 => 0, 2757 => 0, 2758 => 0, 2759 => 0, 2760 => 0, 2761 => 0, 2762 => 0, 2763 => 0, 
2764 => 0, 2765 => 0, 2766 => 0, 2767 => 0, 2768 => 0, 2769 => 0, 2770 => 0, 2771 => 0, 2772 => 0, 2773 => 1, 2774 => 1, 2775 => 1, 2776 => 1, 2777 => 
1, 2778 => 1, 2779 => 1, 2780 => 1, 2781 => 1, 2782 => 1, 2783 => 1, 2784 => 0, 2785 => 0, 2786 => 0, 2787 => 0, 2788 => 0, 2789 => 0, 2790 => 0, 2791 
=> 0, 2792 => 0, 2793 => 0, 2794 => 0, 2795 => 0, 2796 => 0, 2797 => 0, 2798 => 0, 2799 => 0, 2800 => 0, 2801 => 0, 2802 => 0, 2803 => 0, 2804 => 0, 2805 => 1, 2806 => 1, 2807 => 1, 2808 => 1, 2809 => 1, 2810 => 1, 2811 => 1, 2812 => 1, 2813 => 1, 2814 => 1, 2815 => 1, 2816 => 0, 2817 => 0, 2818 => 0, 2819 => 0, 2820 => 0, 2821 => 0, 2822 => 0, 2823 => 0, 2824 => 1, 2825 => 1, 2826 => 1, 2827 => 1, 2828 => 1, 2829 => 1, 2830 => 1, 2831 => 1, 2832 => 1, 2833 => 1, 2834 => 1, 2835 => 0, 2836 => 0, 2837 => 0, 2838 => 0, 2839 => 0, 2840 => 0, 2841 => 0, 2842 => 0, 2843 => 0, 2844 => 0, 2845 => 0, 2846 => 0, 2847 => 0, 2848 => 0, 2849 => 0, 2850 => 0, 2851 => 0, 2852 => 0, 2853 => 0, 2854 => 0, 2855 => 0, 2856 => 1, 2857 => 1, 2858 => 1, 2859 => 1, 2860 => 1, 2861 => 1, 2862 => 1, 2863 => 1, 2864 => 1, 2865 => 1, 2866 => 1, 2867 => 0, 2868 => 0, 2869 => 0, 2870 => 0, 2871 => 0, 2872 => 0, 2873 => 0, 2874 => 0, 2875 => 1, 2876 => 1, 2877 => 1, 2878 => 1, 2879 => 1, 2880 => 1, 2881 => 1, 2882 => 1, 2883 => 1, 2884 => 1, 2885 => 1, 2886 => 1, 2887 => 1, 2888 => 1, 2889 => 1, 2890 => 1, 2891 => 1, 2892 => 1, 2893 => 0, 2894 => 0, 2895 => 0, 2896 => 0, 2897 => 0, 2898 => 0, 2899 => 0, 2900 => 0, 2901 => 0, 2902 => 0, 2903 => 0, 2904 => 0, 2905 => 0, 2906 => 0, 2907 => 1, 2908 => 1, 2909 => 1, 2910 => 1, 2911 => 1, 2912 => 1, 2913 => 1, 2914 => 1, 
2915 => 1, 2916 => 1, 2917 => 1, 2918 => 0, 2919 => 0, 2920 => 0, 2921 => 0, 2922 => 0, 2923 => 0, 2924 => 0, 2925 => 0, 2926 => 1, 2927 => 1, 2928 => 
1, 2929 => 1, 2930 => 1, 2931 => 1, 2932 => 1, 2933 => 1, 2934 => 1, 2935 => 1, 2936 => 1, 2937 => 0, 2938 => 0, 2939 => 0, 2940 => 0, 2941 => 0, 2942 
=> 0, 2943 => 0, 2944 => 0, 2945 => 0, 2946 => 0, 2947 => 0, 2948 => 0, 2949 => 0, 2950 => 0, 2951 => 0, 2952 => 0, 2953 => 0, 2954 => 0, 2955 => 0, 2956 => 0, 2957 => 0, 2958 => 0, 2959 => 0, 2960 => 0, 2961 => 0, 2962 => 0, 2963 => 0, 2964 => 0, 2965 => 0, 2966 => 0, 2967 => 0, 2968 => 0, 2969 => 0, 2970 => 0, 2971 => 1, 2972 => 1, 2973 => 1, 2974 => 1, 2975 => 1, 2976 => 1, 2977 => 1, 2978 => 1, 2979 => 1, 2980 => 1, 2981 => 1, 2982 => 0, 2983 => 0, 2984 => 0, 2985 => 0, 2986 => 0, 2987 => 0, 2988 => 0, 2989 => 0, 2990 => 0, 2991 => 0, 2992 => 0, 2993 => 0, 2994 => 0, 2995 => 0, 2996 => 0, 2997 => 0, 2998 => 0, 2999 => 0, 3000 => 0, 3001 => 0, 3002 => 0, 3003 => 1, 3004 => 1, 3005 => 1, 3006 => 1, 3007 => 1, 3008 => 1, 3009 => 1, 3010 => 1, 3011 => 1, 3012 => 1, 3013 => 1, 3014 => 0, 3015 => 0, 3016 => 0, 3017 => 0, 3018 => 0, 3019 => 0, 3020 => 0, 3021 => 0, 3022 => 1, 3023 => 1, 3024 => 1, 3025 => 1, 3026 => 1, 3027 => 1, 3028 => 1, 3029 => 1, 3030 => 1, 3031 => 1, 3032 => 1, 3033 => 0, 3034 => 0, 3035 => 0, 3036 => 0, 3037 => 0, 3038 => 0, 3039 => 0, 3040 => 0, 3041 => 0, 3042 => 0, 3043 => 0, 3044 => 0, 3045 => 0, 3046 => 0, 3047 => 0, 3048 => 0, 3049 => 0, 3050 => 0, 3051 => 0, 3052 => 0, 3053 => 0, 3054 => 1, 3055 => 1, 3056 => 1, 3057 => 1, 3058 => 1, 3059 => 1, 3060 => 1, 3061 => 1, 3062 => 1, 3063 => 1, 3064 => 1, 3065 => 0, 
3066 => 0, 3067 => 0, 3068 => 0, 3069 => 0, 3070 => 0, 3071 => 0, 3072 => 0, 3073 => 1, 3074 => 1, 3075 => 1, 3076 => 1, 3077 => 1, 3078 => 1, 3079 => 
1, 3080 => 1, 3081 => 1, 3082 => 1, 3083 => 1, 3084 => 1, 3085 => 1, 3086 => 1, 3087 => 1, 3088 => 1, 3089 => 1, 3090 => 1, 3091 => 0, 3092 => 0, 3093 
=> 0, 3094 => 0, 3095 => 0, 3096 => 0, 3097 => 0, 3098 => 0, 3099 => 0, 3100 => 0, 3101 => 0, 3102 => 0, 3103 => 0, 3104 => 0, 3105 => 1, 3106 => 1, 3107 => 1, 3108 => 1, 3109 => 1, 3110 => 1, 3111 => 1, 3112 => 1, 3113 => 1, 3114 => 1, 3115 => 1, 3116 => 0, 3117 => 0, 3118 => 0, 3119 => 0, 3120 => 0, 3121 => 0, 3122 => 0, 3123 => 0, 3124 => 1, 3125 => 1, 3126 => 1, 3127 => 1, 3128 => 1, 3129 => 1, 3130 => 1, 3131 => 1, 3132 => 1, 3133 => 1, 3134 => 1, 3135 => 0, 3136 => 0, 3137 => 0, 3138 => 0, 3139 => 0, 3140 => 0, 3141 => 0, 3142 => 0, 3143 => 0, 3144 => 0, 3145 => 0, 3146 => 0, 3147 => 0, 3148 => 0, 3149 => 0, 3150 => 0, 3151 => 0, 3152 => 0, 3153 => 0, 3154 => 0, 3155 => 0, 3156 => 0, 3157 => 0, 3158 => 0, 3159 => 0, 3160 => 0, 3161 => 0, 3162 => 0, 3163 => 0, 3164 => 0, 3165 => 0, 3166 => 0, 3167 => 0, 3168 => 0, 3169 => 1, 3170 => 1, 3171 => 1, 3172 => 1, 3173 => 1, 3174 => 1, 3175 => 1, 3176 => 1, 3177 => 1, 3178 => 1, 3179 => 1, 3180 => 0, 3181 => 0, 3182 => 0, 3183 => 0, 3184 => 0, 3185 => 0, 3186 => 0, 3187 => 0, 3188 => 0, 3189 => 0, 3190 => 0, 3191 => 0, 3192 => 0, 3193 => 0, 3194 => 0, 3195 => 0, 3196 => 0, 3197 => 0, 3198 => 0, 3199 => 0, 3200 => 0, 3201 => 1, 3202 => 1, 3203 => 1, 3204 => 1, 3205 => 1, 3206 => 1, 3207 => 1, 3208 => 1, 3209 => 1, 3210 => 1, 3211 => 1, 3212 => 0, 3213 => 0, 3214 => 0, 3215 => 0, 3216 => 0, 
3217 => 0, 3218 => 0, 3219 => 0, 3220 => 1, 3221 => 1, 3222 => 1, 3223 => 1, 3224 => 1, 3225 => 1, 3226 => 1, 3227 => 1, 3228 => 1, 3229 => 1, 3230 => 
1, 3231 => 0, 3232 => 0, 3233 => 0, 3234 => 0, 3235 => 0, 3236 => 0, 3237 => 0, 3238 => 0, 3239 => 0, 3240 => 0, 3241 => 0, 3242 => 0, 3243 => 0, 3244 
=> 0, 3245 => 0, 3246 => 0, 3247 => 0, 3248 => 0, 3249 => 0, 3250 => 0, 3251 => 0, 3252 => 1, 3253 => 1, 3254 => 1, 3255 => 1, 3256 => 1, 3257 => 1, 3258 => 1, 3259 => 1, 3260 => 1, 3261 => 1, 3262 => 1, 3263 => 0, 3264 => 0, 3265 => 0, 3266 => 0, 3267 => 0, 3268 => 0, 3269 => 0, 3270 => 0, 3271 => 1, 3272 => 1, 3273 => 1, 3274 => 1, 3275 => 1, 3276 => 1, 3277 => 1, 3278 => 1, 3279 => 1, 3280 => 1, 3281 => 1, 3282 => 1, 3283 => 1, 3284 => 1, 3285 => 1, 3286 => 1, 3287 => 1, 3288 => 1, 3289 => 0, 3290 => 0, 3291 => 0, 3292 => 0, 3293 => 0, 3294 => 0, 3295 => 0, 3296 => 0, 3297 => 0, 3298 => 0, 3299 => 0, 3300 => 0, 3301 => 0, 3302 => 0, 3303 => 1, 3304 => 1, 3305 => 1, 3306 => 1, 3307 => 1, 3308 => 1, 3309 => 1, 3310 => 1, 3311 => 1, 3312 => 1, 3313 => 1, 3314 => 0, 3315 => 0, 3316 => 0, 3317 => 0, 3318 => 0, 3319 => 0, 3320 => 0, 3321 => 0, 3322 => 1, 3323 => 1, 3324 => 1, 3325 => 1, 3326 => 1, 3327 => 1, 3328 => 1, 3329 => 1, 3330 => 1, 3331 => 1, 3332 => 1, 3333 => 0, 3334 => 0, 3335 => 0, 3336 => 0, 3337 => 0, 3338 => 0, 3339 => 0, 3340 => 0, 3341 => 0, 3342 => 0, 3343 => 0, 3344 => 0, 3345 => 0, 3346 => 0, 3347 => 0, 3348 => 0, 3349 => 0, 3350 => 0, 3351 => 0, 3352 => 0, 3353 => 0, 3354 => 0, 3355 => 0, 3356 => 0, 3357 => 0, 3358 => 0, 3359 => 0, 3360 => 0, 3361 => 0, 3362 => 0, 3363 => 0, 3364 => 0, 3365 => 0, 3366 => 0, 3367 => 1, 
3368 => 1, 3369 => 1, 3370 => 1, 3371 => 1, 3372 => 1, 3373 => 1, 3374 => 1, 3375 => 1, 3376 => 1, 3377 => 1, 3378 => 0, 3379 => 0, 3380 => 0, 3381 => 
0, 3382 => 0, 3383 => 0, 3384 => 0, 3385 => 0, 3386 => 0, 3387 => 0, 3388 => 0, 3389 => 0, 3390 => 0, 3391 => 0, 3392 => 0, 3393 => 0, 3394 => 0, 3395 
=> 0, 3396 => 0, 3397 => 0, 3398 => 0, 3399 => 1, 3400 => 1, 3401 => 1, 3402 => 1, 3403 => 1, 3404 => 1, 3405 => 1, 3406 => 1, 3407 => 1, 3408 => 1, 3409 => 1, 3410 => 0, 3411 => 0, 3412 => 0, 3413 => 0, 3414 => 0, 3415 => 0, 3416 => 0, 3417 => 0, 3418 => 1, 3419 => 1, 3420 => 1, 3421 => 1, 3422 => 1, 3423 => 1, 3424 => 1, 3425 => 1, 3426 => 1, 3427 => 1, 3428 => 1, 3429 => 0, 3430 => 0, 3431 => 0, 3432 => 0, 3433 => 0, 3434 => 0, 3435 => 0, 3436 => 0, 3437 => 0, 3438 => 0, 3439 => 0, 3440 => 0, 3441 => 0, 3442 => 0, 3443 => 0, 3444 => 0, 3445 => 0, 3446 => 0, 3447 => 0, 3448 => 0, 3449 => 0, 3450 => 1, 3451 => 1, 3452 => 1, 3453 => 1, 3454 => 1, 3455 => 1, 3456 => 1, 3457 => 1, 3458 => 1, 3459 => 1, 3460 => 1, 3461 => 0, 3462 => 0, 3463 => 0, 3464 => 0, 3465 => 0, 3466 => 0, 3467 => 0, 3468 => 0, 3469 => 1, 3470 => 1, 3471 => 1, 3472 => 1, 3473 => 1, 3474 => 1, 3475 => 1, 3476 => 1, 3477 => 1, 3478 => 1, 3479 => 1, 3480 => 1, 3481 => 1, 3482 => 1, 3483 => 1, 3484 => 1, 3485 => 1, 3486 => 1, 3487 => 0, 3488 => 0, 3489 => 0, 3490 => 0, 3491 => 0, 3492 => 0, 3493 => 0, 3494 => 0, 3495 => 0, 3496 => 0, 3497 => 0, 3498 => 0, 3499 => 0, 3500 => 0, 3501 => 1, 3502 => 1, 3503 => 1, 3504 => 1, 3505 => 1, 3506 => 1, 3507 => 1, 3508 => 1, 3509 => 1, 3510 => 1, 3511 => 1, 3512 => 0, 3513 => 0, 3514 => 0, 3515 => 0, 3516 => 0, 3517 => 0, 3518 => 0, 
3519 => 0, 3520 => 1, 3521 => 1, 3522 => 1, 3523 => 1, 3524 => 1, 3525 => 1, 3526 => 1, 3527 => 1, 3528 => 1, 3529 => 1, 3530 => 1, 3531 => 0, 3532 => 
0, 3533 => 0, 3534 => 0, 3535 => 0, 3536 => 0, 3537 => 0, 3538 => 0, 3539 => 0, 3540 => 0, 3541 => 0, 3542 => 0, 3543 => 0, 3544 => 0, 3545 => 0, 3546 
=> 0, 3547 => 0, 3548 => 0, 3549 => 0, 3550 => 0, 3551 => 0, 3552 => 0, 3553 => 0, 3554 => 0, 3555 => 0, 3556 => 0, 3557 => 0, 3558 => 0, 3559 => 0, 3560 => 0, 3561 => 0, 3562 => 0, 3563 => 0, 3564 => 0, 3565 => 1, 3566 => 1, 3567 => 1, 3568 => 1, 3569 => 1, 3570 => 1, 3571 => 1, 3572 => 1, 3573 => 1, 3574 => 1, 3575 => 1, 3576 => 0, 3577 => 0, 3578 => 0, 3579 => 0, 3580 => 0, 3581 => 0, 3582 => 0, 3583 => 0, 3584 => 0, 3585 => 0, 3586 => 0, 3587 => 0, 3588 => 0, 3589 => 0, 3590 => 0, 3591 => 0, 3592 => 0, 3593 => 0, 3594 => 0, 3595 => 0, 3596 => 0, 3597 => 1, 3598 => 1, 3599 => 1, 3600 => 1, 3601 => 1, 3602 => 1, 3603 => 1, 3604 => 1, 3605 => 1, 3606 => 1, 3607 => 1, 3608 => 0, 3609 => 0, 3610 => 0, 3611 => 0, 3612 => 0, 3613 => 0, 3614 => 0, 3615 => 0, 3616 => 1, 3617 => 1, 3618 => 1, 3619 => 1, 3620 => 1, 3621 => 1, 3622 => 1, 3623 => 1, 3624 => 1, 3625 => 1, 3626 => 1, 3627 => 0, 3628 => 0, 3629 => 0, 3630 => 0, 3631 => 0, 3632 => 0, 3633 => 0, 3634 => 0, 3635 => 0, 3636 => 0, 3637 => 0, 3638 => 0, 3639 => 0, 3640 => 0, 3641 => 0, 3642 => 0, 3643 => 0, 3644 => 0, 3645 => 0, 3646 => 0, 3647 => 0, 3648 => 1, 3649 => 1, 3650 => 1, 3651 => 1, 3652 => 1, 3653 => 1, 3654 => 1, 3655 => 1, 3656 => 1, 3657 => 1, 3658 => 1, 3659 => 0, 3660 => 0, 3661 => 0, 3662 => 0, 3663 => 0, 3664 => 0, 3665 => 0, 3666 => 0, 3667 => 1, 3668 => 1, 3669 => 1, 
3670 => 1, 3671 => 1, 3672 => 1, 3673 => 1, 3674 => 1, 3675 => 1, 3676 => 1, 3677 => 1, 3678 => 1, 3679 => 1, 3680 => 1, 3681 => 1, 3682 => 1, 3683 => 
1, 3684 => 1, 3685 => 0, 3686 => 0, 3687 => 0, 3688 => 0, 3689 => 0, 3690 => 0, 3691 => 0, 3692 => 0, 3693 => 0, 3694 => 0, 3695 => 0, 3696 => 0, 3697 
=> 0, 3698 => 0, 3699 => 1, 3700 => 1, 3701 => 1, 3702 => 1, 3703 => 1, 3704 => 1, 3705 => 1, 3706 => 1, 3707 => 1, 3708 => 1, 3709 => 1, 3710 => 0, 3711 => 0, 3712 => 0, 3713 => 0, 3714 => 0, 3715 => 0, 3716 => 0, 3717 => 0, 3718 => 1, 3719 => 1, 3720 => 1, 3721 => 1, 3722 => 1, 3723 => 1, 3724 => 1, 3725 => 1, 3726 => 1, 3727 => 1, 3728 => 1, 3729 => 0, 3730 => 0, 3731 => 0, 3732 => 0, 3733 => 0, 3734 => 0, 3735 => 0, 3736 => 0, 3737 => 0, 3738 => 0, 3739 => 0, 3740 => 0, 3741 => 0, 3742 => 0, 3743 => 0, 3744 => 0, 3745 => 0, 3746 => 0, 3747 => 0, 3748 => 0, 3749 => 0, 3750 => 0, 3751 => 0, 3752 => 0, 3753 => 0, 3754 => 0, 3755 => 0, 3756 => 0, 3757 => 0, 3758 => 0, 3759 => 0, 3760 => 0, 3761 => 0, 3762 => 0, 3763 => 1, 3764 => 1, 3765 => 1, 3766 => 1, 3767 => 1, 3768 => 1, 3769 => 1, 3770 => 1, 3771 => 1, 3772 => 1, 3773 => 1, 3774 => 0, 3775 => 0, 3776 => 0, 3777 => 0, 3778 => 0, 3779 => 0, 3780 => 0, 3781 => 0, 3782 => 0, 3783 => 0, 3784 => 0, 3785 => 0, 3786 => 0, 3787 => 0, 3788 => 0, 3789 => 0, 3790 => 0, 3791 => 0, 3792 => 0, 3793 => 0, 3794 => 0, 3795 => 1, 3796 => 1, 3797 => 1, 3798 => 1, 3799 => 1, 3800 => 1, 3801 => 1, 3802 => 1, 3803 => 1, 3804 => 1, 3805 => 1, 3806 => 0, 3807 => 0, 3808 => 0, 3809 => 0, 3810 => 0, 3811 => 0, 3812 => 0, 3813 => 0, 3814 => 1, 3815 => 1, 3816 => 1, 3817 => 1, 3818 => 1, 3819 => 1, 3820 => 1, 
3821 => 1, 3822 => 1, 3823 => 1, 3824 => 1, 3825 => 0, 3826 => 0, 3827 => 0, 3828 => 0, 3829 => 0, 3830 => 0, 3831 => 0, 3832 => 0, 3833 => 0, 3834 => 
0, 3835 => 0, 3836 => 0, 3837 => 0, 3838 => 0, 3839 => 0, 3840 => 0, 3841 => 0, 3842 => 0, 3843 => 0, 3844 => 0, 3845 => 0, 3846 => 1, 3847 => 1, 3848 
=> 1, 3849 => 1, 3850 => 1, 3851 => 1, 3852 => 1, 3853 => 1, 3854 => 1, 3855 => 1, 3856 => 1, 3857 => 0, 3858 => 0, 3859 => 0, 3860 => 0, 3861 => 0, 3862 => 0, 3863 => 0, 3864 => 0, 3865 => 1, 3866 => 1, 3867 => 1, 3868 => 1, 3869 => 1, 3870 => 1, 3871 => 1, 3872 => 1, 3873 => 1, 3874 => 1, 3875 => 1, 3876 => 0, 3877 => 0, 3878 => 0, 3879 => 0, 3880 => 0, 3881 => 0, 3882 => 0, 3883 => 0, 3884 => 0, 3885 => 0, 3886 => 0, 3887 => 0, 3888 => 0, 3889 => 0, 3890 => 0, 3891 => 0, 3892 => 0, 3893 => 0, 3894 => 0, 3895 => 0, 3896 => 0, 3897 => 1, 3898 => 1, 3899 => 1, 3900 => 1, 3901 => 1, 3902 => 1, 3903 => 1, 3904 => 1, 3905 => 1, 3906 => 1, 3907 => 1, 3908 => 0, 3909 => 0, 3910 => 0, 3911 => 0, 3912 => 0, 3913 => 0, 3914 => 0, 3915 => 0, 3916 => 1, 3917 => 1, 3918 => 1, 3919 => 1, 3920 => 1, 3921 => 1, 3922 => 1, 3923 => 1, 3924 => 1, 3925 => 1, 3926 => 1, 3927 => 0, 3928 => 0, 3929 => 0, 3930 => 0, 3931 => 0, 3932 => 0, 3933 => 0, 3934 => 0, 3935 => 0, 3936 => 0, 3937 => 0, 3938 => 0, 3939 => 0, 3940 => 0, 3941 => 0, 3942 => 0, 3943 => 0, 3944 => 0, 3945 => 0, 3946 => 0, 3947 => 0, 3948 => 0, 3949 => 0, 3950 => 0, 3951 => 0, 3952 => 0, 3953 => 0, 3954 => 0, 3955 => 0, 3956 => 0, 3957 => 0, 3958 => 0, 3959 => 0, 3960 => 0, 3961 => 1, 3962 => 1, 3963 => 1, 3964 => 1, 3965 => 1, 3966 => 1, 3967 => 1, 3968 => 1, 3969 => 1, 3970 => 1, 3971 => 1, 
3972 => 0, 3973 => 0, 3974 => 0, 3975 => 0, 3976 => 0, 3977 => 0, 3978 => 0, 3979 => 0, 3980 => 0, 3981 => 0, 3982 => 0, 3983 => 0, 3984 => 0, 3985 => 
0, 3986 => 0, 3987 => 0, 3988 => 0, 3989 => 0, 3990 => 0, 3991 => 0, 3992 => 0, 3993 => 1, 3994 => 1, 3995 => 1, 3996 => 1, 3997 => 1, 3998 => 1, 3999 
=> 1, 4000 => 1, 4001 => 1, 4002 => 1, 4003 => 1, 4004 => 0, 4005 => 0, 4006 => 0, 4007 => 0, 4008 => 0, 4009 => 0, 4010 => 0, 4011 => 0, 4012 => 1, 4013 => 1, 4014 => 1, 4015 => 1, 4016 => 1, 4017 => 1, 4018 => 1, 4019 => 1, 4020 => 1, 4021 => 1, 4022 => 1, 4023 => 0, 4024 => 0, 4025 => 0, 4026 => 0, 4027 => 0, 4028 => 0, 4029 => 0, 4030 => 0, 4031 => 0, 4032 => 0, 4033 => 0, 4034 => 0, 4035 => 0, 4036 => 0, 4037 => 0, 4038 => 0, 4039 => 0, 4040 => 0, 4041 => 0, 4042 => 0, 4043 => 0, 4044 => 1, 4045 => 1, 4046 => 1, 4047 => 1, 4048 => 1, 4049 => 1, 4050 => 1, 4051 => 1, 4052 => 1, 4053 => 1, 4054 => 1, 4055 => 0, 4056 => 0, 4057 => 0, 4058 => 0, 4059 => 0, 4060 => 0, 4061 => 0, 4062 => 0, 4063 => 1, 4064 => 1, 4065 => 1, 4066 => 1, 4067 => 1, 4068 => 1, 4069 => 1, 4070 => 1, 4071 => 1, 4072 => 1, 4073 => 1, 4074 => 0, 4075 => 0, 4076 => 0, 4077 => 0, 4078 => 0, 4079 => 0, 4080 => 0, 4081 => 0, 4082 => 1, 4083 => 1, 4084 => 1, 4085 => 1, 4086 => 1, 4087 => 0, 4088 => 0, 4089 => 0, 4090 => 0, 4091 => 0, 4092 => 0, 4093 => 0, 4094 => 0, 4095 => 1, 4096 => 1, 4097 => 1, 4098 => 1, 4099 => 1, 4100 => 1, 4101 => 1, 4102 => 1, 4103 => 1, 4104 => 1, 4105 => 1, 4106 => 0, 4107 => 0, 4108 => 0, 4109 => 0, 4110 => 0, 4111 => 0, 4112 => 0, 4113 => 0, 4114 => 1, 4115 => 1, 4116 => 1, 4117 => 1, 4118 => 1, 4119 => 1, 4120 => 1, 4121 => 1, 4122 => 1, 
4123 => 1, 4124 => 1, 4125 => 0, 4126 => 0, 4127 => 0, 4128 => 0, 4129 => 0, 4130 => 0, 4131 => 0, 4132 => 0, 4133 => 1, 4134 => 1, 4135 => 1, 4136 => 
1, 4137 => 1, 4138 => 1, 4139 => 1, 4140 => 1, 4141 => 1, 4142 => 1, 4143 => 1, 4144 => 1, 4145 => 1, 4146 => 1, 4147 => 1, 4148 => 1, 4149 => 1, 4150 
=> 1, 4151 => 1, 4152 => 1, 4153 => 1, 4154 => 1, 4155 => 1, 4156 => 1, 4157 => 0, 4158 => 0, 4159 => 1, 4160 => 1, 4161 => 1, 4162 => 1, 4163 => 1, 4164 => 1, 4165 => 1, 4166 => 1, 4167 => 1, 4168 => 1, 4169 => 1, 4170 => 0, 4171 => 0, 4172 => 0, 4173 => 0, 4174 => 0, 4175 => 0, 4176 => 0, 4177 => 0, 4178 => 0, 4179 => 0, 4180 => 0, 4181 => 0, 4182 => 0, 4183 => 0, 4184 => 0, 4185 => 0, 4186 => 0, 4187 => 0, 4188 => 0, 4189 => 0, 4190 => 0, 4191 => 1, 4192 => 1, 4193 => 1, 4194 => 1, 4195 => 1, 4196 => 1, 4197 => 1, 4198 => 1, 4199 => 1, 4200 => 1, 4201 => 1, 4202 => 0, 4203 => 0, 4204 => 0, 4205 => 0, 4206 => 0, 4207 => 0, 4208 => 0, 4209 => 0, 4210 => 1, 4211 => 1, 4212 => 1, 4213 => 1, 4214 => 1, 4215 => 1, 4216 => 1, 4217 => 1, 4218 => 1, 4219 => 1, 4220 => 1, 4221 => 0, 4222 => 0, 4223 => 0, 4224 => 0, 4225 => 0, 4226 => 0, 4227 => 0, 4228 => 0, 4229 => 0, 4230 => 0, 4231 => 0, 4232 => 0, 4233 => 0, 4234 => 0, 4235 => 0, 4236 => 0, 4237 => 0, 4238 => 0, 4239 => 0, 4240 => 0, 4241 => 0, 4242 => 1, 4243 => 1, 4244 => 1, 4245 => 1, 4246 => 1, 4247 => 1, 4248 => 1, 4249 => 1, 4250 => 1, 4251 => 1, 4252 => 1, 4253 => 0, 4254 => 0, 4255 => 0, 4256 => 0, 4257 => 0, 4258 => 0, 4259 => 0, 4260 => 0, 4261 => 1, 4262 => 1, 4263 => 1, 4264 => 1, 4265 => 1, 4266 => 1, 4267 => 1, 4268 => 1, 4269 => 1, 4270 => 1, 4271 => 1, 4272 => 0, 4273 => 0, 
4274 => 0, 4275 => 0, 4276 => 0, 4277 => 0, 4278 => 0, 4279 => 0, 4280 => 1, 4281 => 1, 4282 => 1, 4283 => 1, 4284 => 1, 4285 => 0, 4286 => 0, 4287 => 
0, 4288 => 0, 4289 => 0, 4290 => 0, 4291 => 0, 4292 => 0, 4293 => 1, 4294 => 1, 4295 => 1, 4296 => 1, 4297 => 1, 4298 => 1, 4299 => 1, 4300 => 1, 4301 
=> 1, 4302 => 1, 4303 => 1, 4304 => 0, 4305 => 0, 4306 => 0, 4307 => 0, 4308 => 0, 4309 => 0, 4310 => 0, 4311 => 0, 4312 => 1, 4313 => 1, 4314 => 1, 4315 => 1, 4316 => 1, 4317 => 1, 4318 => 1, 4319 => 1, 4320 => 1, 4321 => 1, 4322 => 1, 4323 => 0, 4324 => 0, 4325 => 0, 4326 => 0, 4327 => 0, 4328 => 0, 4329 => 0, 4330 => 0, 4331 => 1, 4332 => 1, 4333 => 1, 4334 => 1, 4335 => 1, 4336 => 1, 4337 => 1, 4338 => 1, 4339 => 1, 4340 => 1, 4341 => 1, 4342 => 1, 4343 => 1, 4344 => 1, 4345 => 1, 4346 => 1, 4347 => 1, 4348 => 1, 4349 => 1, 4350 => 1, 4351 => 1, 4352 => 1, 4353 => 1, 4354 => 1, 4355 => 0, 4356 => 0, 4357 => 1, 4358 => 1, 4359 => 1, 4360 => 1, 4361 => 1, 4362 => 1, 4363 => 1, 4364 => 1, 4365 => 1, 4366 => 1, 4367 => 1, 4368 => 0, 4369 => 0, 4370 => 0, 4371 => 0, 4372 => 0, 4373 => 0, 4374 => 0, 4375 => 0, 4376 => 0, 4377 => 0, 4378 => 0, 4379 => 0, 4380 => 0, 4381 => 0, 4382 => 0, 4383 => 0, 4384 => 0, 4385 => 0, 4386 => 0, 4387 => 0, 4388 => 0, 4389 => 1, 4390 => 1, 4391 => 1, 4392 => 1, 4393 => 1, 4394 => 1, 4395 => 1, 4396 => 1, 4397 => 1, 4398 => 1, 4399 => 1, 4400 => 0, 4401 => 0, 4402 => 0, 4403 => 0, 4404 => 0, 4405 => 0, 4406 => 0, 4407 => 0, 4408 => 1, 4409 => 1, 4410 => 1, 4411 => 1, 4412 => 1, 4413 => 1, 4414 => 1, 4415 => 1, 4416 => 1, 4417 => 1, 4418 => 1, 4419 => 0, 4420 => 0, 4421 => 0, 4422 => 0, 4423 => 0, 4424 => 0, 
4425 => 0, 4426 => 0, 4427 => 0, 4428 => 0, 4429 => 0, 4430 => 0, 4431 => 0, 4432 => 0, 4433 => 0, 4434 => 0, 4435 => 0, 4436 => 0, 4437 => 0, 4438 => 
0, 4439 => 0, 4440 => 1, 4441 => 1, 4442 => 1, 4443 => 1, 4444 => 1, 4445 => 1, 4446 => 1, 4447 => 1, 4448 => 1, 4449 => 1, 4450 => 1, 4451 => 0, 4452 
=> 0, 4453 => 0, 4454 => 0, 4455 => 0, 4456 => 0, 4457 => 0, 4458 => 0, 4459 => 1, 4460 => 1, 4461 => 1, 4462 => 1, 4463 => 1, 4464 => 1, 4465 => 1, 4466 => 1, 4467 => 1, 4468 => 1, 4469 => 1, 4470 => 0, 4471 => 0, 4472 => 0, 4473 => 0, 4474 => 0, 4475 => 0, 4476 => 0, 4477 => 0, 4478 => 1, 4479 => 1, 4480 => 1, 4481 => 1, 4482 => 1, 4483 => 0, 4484 => 0, 4485 => 0, 4486 => 0, 4487 => 0, 4488 => 0, 4489 => 0, 4490 => 0, 4491 => 1, 4492 => 1, 4493 => 1, 4494 => 1, 4495 => 1, 4496 => 1, 4497 => 1, 4498 => 1, 4499 => 1, 4500 => 1, 4501 => 1, 4502 => 0, 4503 => 0, 4504 => 0, 4505 => 0, 4506 => 0, 4507 => 0, 4508 => 0, 4509 => 0, 4510 => 1, 4511 => 1, 4512 => 1, 4513 => 1, 4514 => 1, 4515 => 1, 4516 => 1, 4517 => 1, 4518 => 1, 4519 => 1, 4520 => 1, 4521 => 0, 4522 => 0, 4523 => 0, 4524 => 0, 4525 => 0, 4526 => 0, 4527 => 0, 4528 => 0, 4529 => 1, 4530 => 1, 4531 => 1, 4532 => 1, 4533 => 1, 4534 => 1, 4535 => 1, 4536 => 1, 4537 => 1, 4538 => 1, 4539 => 1, 4540 => 1, 4541 => 1, 4542 => 1, 4543 => 1, 4544 => 1, 4545 => 1, 4546 => 1, 4547 => 1, 4548 => 1, 4549 => 1, 4550 => 1, 4551 => 1, 4552 => 1, 4553 => 0, 4554 => 0, 4555 => 1, 4556 => 1, 4557 => 1, 4558 => 1, 4559 => 1, 4560 => 1, 4561 => 1, 4562 => 1, 4563 => 1, 4564 => 1, 4565 => 1, 4566 => 0, 4567 => 0, 4568 => 0, 4569 => 0, 4570 => 0, 4571 => 0, 4572 => 0, 4573 => 0, 4574 => 0, 4575 => 0, 
4576 => 0, 4577 => 0, 4578 => 0, 4579 => 0, 4580 => 0, 4581 => 0, 4582 => 0, 4583 => 0, 4584 => 0, 4585 => 0, 4586 => 0, 4587 => 1, 4588 => 1, 4589 => 
1, 4590 => 1, 4591 => 1, 4592 => 1, 4593 => 1, 4594 => 1, 4595 => 1, 4596 => 1, 4597 => 1, 4598 => 0, 4599 => 0, 4600 => 0, 4601 => 0, 4602 => 0, 4603 
=> 0, 4604 => 0, 4605 => 0, 4606 => 1, 4607 => 1, 4608 => 1, 4609 => 1, 4610 => 1, 4611 => 1, 4612 => 1, 4613 => 1, 4614 => 1, 4615 => 1, 4616 => 1, 4617 => 0, 4618 => 0, 4619 => 0, 4620 => 0, 4621 => 0, 4622 => 0, 4623 => 0, 4624 => 0, 4625 => 0, 4626 => 0, 4627 => 0, 4628 => 0, 4629 => 0, 4630 => 0, 4631 => 0, 4632 => 0, 4633 => 0, 4634 => 0, 4635 => 0, 4636 => 0, 4637 => 0, 4638 => 1, 4639 => 1, 4640 => 1, 4641 => 1, 4642 => 1, 4643 => 1, 4644 => 1, 4645 => 1, 4646 => 1, 4647 => 1, 4648 => 1, 4649 => 0, 4650 => 0, 4651 => 0, 4652 => 0, 4653 => 0, 4654 => 0, 4655 => 0, 4656 => 0, 4657 => 1, 4658 => 1, 4659 => 1, 4660 => 1, 4661 => 1, 4662 => 1, 4663 => 1, 4664 => 1, 4665 => 1, 4666 => 1, 4667 => 1, 4668 => 0, 4669 => 0, 4670 => 0, 4671 => 0, 4672 => 0, 4673 => 0, 4674 => 0, 4675 => 0, 4676 => 1, 4677 => 1, 4678 => 1, 4679 => 1, 4680 => 1, 4681 => 0, 4682 => 0, 4683 => 0, 4684 => 0, 4685 => 0, 4686 => 0, 4687 => 0, 4688 => 0, 4689 => 1, 4690 => 1, 4691 => 1, 4692 => 1, 4693 => 1, 4694 => 1, 4695 => 1, 4696 => 1, 4697 => 1, 4698 => 1, 4699 => 1, 4700 => 0, 4701 => 0, 4702 => 0, 4703 => 0, 4704 => 0, 4705 => 0, 4706 => 0, 4707 => 0, 4708 => 1, 4709 => 1, 4710 => 1, 4711 => 1, 4712 => 1, 4713 => 1, 4714 => 1, 4715 => 1, 4716 => 1, 4717 => 1, 4718 => 1, 4719 => 0, 4720 => 0, 4721 => 0, 4722 => 0, 4723 => 0, 4724 => 0, 4725 => 0, 4726 => 0, 
4727 => 1, 4728 => 1, 4729 => 1, 4730 => 1, 4731 => 1, 4732 => 1, 4733 => 1, 4734 => 1, 4735 => 1, 4736 => 1, 4737 => 1, 4738 => 1, 4739 => 1, 4740 => 
1, 4741 => 1, 4742 => 1, 4743 => 1, 4744 => 1, 4745 => 1, 4746 => 1, 4747 => 1, 4748 => 1, 4749 => 1, 4750 => 1, 4751 => 0, 4752 => 0, 4753 => 1, 4754 
=> 1, 4755 => 1, 4756 => 1, 4757 => 1, 4758 => 1, 4759 => 1, 4760 => 1, 4761 => 1, 4762 => 1, 4763 => 1, 4764 => 0, 4765 => 0, 4766 => 0, 4767 => 0, 4768 => 0, 4769 => 0, 4770 => 0, 4771 => 0, 4772 => 0, 4773 => 0, 4774 => 0, 4775 => 0, 4776 => 0, 4777 => 0, 4778 => 0, 4779 => 0, 4780 => 0, 4781 => 0, 4782 => 0, 4783 => 0, 4784 => 0, 4785 => 1, 4786 => 1, 4787 => 1, 4788 => 1, 4789 => 1, 4790 => 1, 4791 => 1, 4792 => 1, 4793 => 1, 4794 => 1, 4795 => 1, 4796 => 0, 4797 => 0, 4798 => 0, 4799 => 0, 4800 => 0, 4801 => 0, 4802 => 0, 4803 => 0, 4804 => 1, 4805 => 1, 4806 => 1, 4807 => 1, 4808 => 1, 4809 => 1, 4810 => 1, 4811 => 1, 4812 => 1, 4813 => 1, 4814 => 1, 4815 => 0, 4816 => 0, 4817 => 0, 4818 => 0, 4819 => 0, 4820 => 0, 4821 => 0, 4822 => 0, 4823 => 0, 4824 => 0, 4825 => 0, 4826 => 0, 4827 => 0, 4828 => 0, 4829 => 0, 4830 => 0, 4831 => 0, 4832 => 0, 4833 => 0, 4834 => 0, 4835 => 0, 4836 => 1, 4837 => 1, 4838 => 1, 4839 => 1, 4840 => 1, 4841 => 1, 4842 => 1, 4843 => 1, 4844 => 1, 4845 => 1, 4846 => 1, 4847 => 0, 4848 => 0, 4849 => 0, 4850 => 0, 4851 => 0, 4852 => 0, 4853 => 0, 4854 => 0, 4855 => 1, 4856 => 1, 4857 => 1, 4858 => 1, 4859 => 1, 4860 => 1, 4861 => 1, 4862 => 1, 4863 => 1, 4864 => 1, 4865 => 1, 4866 => 0, 4867 => 0, 4868 => 0, 4869 => 0, 4870 => 0, 4871 => 0, 4872 => 0, 4873 => 0, 4874 => 1, 4875 => 1, 4876 => 1, 4877 => 1, 
4878 => 1, 4879 => 0, 4880 => 0, 4881 => 0, 4882 => 0, 4883 => 0, 4884 => 0, 4885 => 0, 4886 => 0, 4887 => 1, 4888 => 1, 4889 => 1, 4890 => 1, 4891 => 
1, 4892 => 1, 4893 => 1, 4894 => 1, 4895 => 1, 4896 => 1, 4897 => 1, 4898 => 0, 4899 => 0, 4900 => 0, 4901 => 0, 4902 => 0, 4903 => 0, 4904 => 0, 4905 
=> 0, 4906 => 1, 4907 => 1, 4908 => 1, 4909 => 1, 4910 => 1, 4911 => 1, 4912 => 1, 4913 => 1, 4914 => 1, 4915 => 1, 4916 => 1, 4917 => 0, 4918 => 0, 4919 => 0, 4920 => 0, 4921 => 0, 4922 => 0, 4923 => 0, 4924 => 0, 4925 => 1, 4926 => 1, 4927 => 1, 4928 => 1, 4929 => 1, 4930 => 1, 4931 => 1, 4932 => 1, 4933 => 1, 4934 => 1, 4935 => 1, 4936 => 1, 4937 => 1, 4938 => 1, 4939 => 1, 4940 => 1, 4941 => 1, 4942 => 1, 4943 => 1, 4944 => 1, 4945 => 1, 4946 => 1, 4947 => 1, 4948 => 1, 4949 => 0, 4950 => 0, 4951 => 1, 4952 => 1, 4953 => 1, 4954 => 1, 4955 => 1, 4956 => 1, 4957 => 1, 4958 => 1, 4959 => 1, 4960 => 1, 4961 => 1, 4962 => 0, 4963 => 0, 4964 => 0, 4965 => 0, 4966 => 0, 4967 => 0, 4968 => 0, 4969 => 0, 4970 => 0, 4971 => 0, 4972 => 0, 4973 => 0, 4974 => 0, 4975 => 0, 4976 => 0, 4977 => 0, 4978 => 0, 4979 => 0, 4980 => 0, 4981 => 0, 4982 => 0, 4983 => 1, 4984 => 1, 4985 => 1, 4986 => 1, 4987 => 1, 4988 => 0, 4989 => 0, 4990 => 0, 4991 => 0, 4992 => 0, 4993 => 0, 4994 => 0, 4995 => 0, 4996 => 0, 4997 => 0, 4998 => 0, 4999 => 0, 5000 => 0, 5001 => 0, 5002 => 1, 5003 => 1, 5004 => 1, 5005 => 1, 5006 => 1, 5007 => 1, 5008 => 1, 5009 => 1, 5010 => 1, 5011 => 1, 5012 => 1, 5013 => 0, 5014 => 0, 5015 => 0, 5016 => 0, 5017 => 0, 5018 => 0, 5019 => 0, 5020 => 0, 5021 => 0, 5022 => 0, 5023 => 0, 5024 => 0, 5025 => 0, 5026 => 0, 5027 => 0, 5028 => 0, 
5029 => 0, 5030 => 0, 5031 => 0, 5032 => 0, 5033 => 0, 5034 => 1, 5035 => 1, 5036 => 1, 5037 => 1, 5038 => 1, 5039 => 1, 5040 => 1, 5041 => 1, 5042 => 
1, 5043 => 1, 5044 => 1, 5045 => 0, 5046 => 0, 5047 => 0, 5048 => 0, 5049 => 0, 5050 => 0, 5051 => 0, 5052 => 0, 5053 => 1, 5054 => 1, 5055 => 1, 5056 
=> 1, 5057 => 1, 5058 => 1, 5059 => 1, 5060 => 1, 5061 => 1, 5062 => 1, 5063 => 1, 5064 => 0, 5065 => 0, 5066 => 0, 5067 => 0, 5068 => 0, 5069 => 0, 5070 => 0, 5071 => 0, 5072 => 0, 5073 => 0, 5074 => 0, 5075 => 0, 5076 => 0, 5077 => 0, 5078 => 0, 5079 => 0, 5080 => 0, 5081 => 0, 5082 => 0, 5083 => 0, 5084 => 0, 5085 => 1, 5086 => 1, 5087 => 1, 5088 => 1, 5089 => 1, 5090 => 1, 5091 => 1, 5092 => 1, 5093 => 1, 5094 => 1, 5095 => 1, 5096 => 0, 5097 => 0, 5098 => 0, 5099 => 0, 5100 => 0, 5101 => 0, 5102 => 0, 5103 => 0, 5104 => 1, 5105 => 1, 5106 => 1, 5107 => 1, 5108 => 1, 5109 => 1, 5110 => 1, 5111 => 1, 5112 => 1, 5113 => 1, 5114 => 1, 5115 => 0, 5116 => 0, 5117 => 0, 5118 => 0, 5119 => 0, 5120 => 0, 5121 => 0, 5122 => 0, 5123 => 0, 5124 => 0, 5125 => 0, 5126 => 0, 5127 => 0, 5128 => 0, 5129 => 0, 5130 => 0, 5131 => 0, 5132 => 0, 5133 => 0, 5134 => 0, 5135 => 0, 5136 => 1, 5137 => 1, 5138 => 1, 5139 => 1, 5140 => 1, 5141 => 1, 5142 => 1, 5143 => 1, 5144 => 1, 5145 => 1, 5146 => 1, 5147 => 0, 5148 => 0, 5149 => 1, 5150 => 1, 5151 => 1, 5152 => 1, 5153 => 1, 5154 => 1, 5155 => 1, 5156 => 1, 5157 => 1, 5158 => 1, 5159 => 1, 5160 => 1, 5161 => 1, 5162 => 1, 5163 => 1, 5164 => 1, 5165 => 1, 5166 => 1, 5167 => 1, 5168 => 1, 5169 => 1, 5170 => 1, 5171 => 1, 5172 => 1, 5173 => 1, 5174 => 1, 5175 => 1, 5176 => 1, 5177 => 1, 5178 => 1, 5179 => 1, 
5180 => 1, 5181 => 1, 5182 => 1, 5183 => 1, 5184 => 1, 5185 => 0, 5186 => 0, 5187 => 0, 5188 => 0, 5189 => 0, 5190 => 0, 5191 => 0, 5192 => 0, 5193 => 
0, 5194 => 0, 5195 => 0, 5196 => 0, 5197 => 0, 5198 => 0, 5199 => 0, 5200 => 1, 5201 => 1, 5202 => 1, 5203 => 1, 5204 => 1, 5205 => 1, 5206 => 1, 5207 
=> 1, 5208 => 1, 5209 => 1, 5210 => 1, 5211 => 0, 5212 => 0, 5213 => 0, 5214 => 0, 5215 => 0, 5216 => 0, 5217 => 0, 5218 => 0, 5219 => 0, 5220 => 0, 5221 => 0, 5222 => 0, 5223 => 0, 5224 => 0, 5225 => 0, 5226 => 0, 5227 => 0, 5228 => 0, 5229 => 0, 5230 => 0, 5231 => 0, 5232 => 1, 5233 => 1, 5234 => 1, 5235 => 1, 5236 => 1, 5237 => 1, 5238 => 1, 5239 => 1, 5240 => 1, 5241 => 1, 5242 => 1, 5243 => 0, 5244 => 0, 5245 => 0, 5246 => 0, 5247 => 0, 5248 => 0, 5249 => 0, 5250 => 0, 5251 => 1, 5252 => 1, 5253 => 1, 5254 => 1, 5255 => 1, 5256 => 1, 5257 => 1, 5258 => 1, 5259 => 1, 5260 => 1, 5261 => 1, 5262 => 0, 5263 => 0, 5264 => 0, 5265 => 0, 5266 => 0, 5267 => 0, 5268 => 0, 5269 => 0, 5270 => 0, 5271 => 0, 5272 => 0, 5273 => 0, 5274 => 0, 5275 => 0, 5276 => 1, 5277 => 1, 5278 => 1, 5279 => 1, 5280 => 1, 5281 => 1, 5282 => 1, 5283 => 1, 5284 => 1, 5285 => 1, 5286 => 1, 5287 => 1, 5288 => 1, 5289 => 1, 5290 => 1, 5291 => 1, 5292 => 1, 5293 => 1, 5294 => 0, 5295 => 0, 5296 => 0, 5297 => 0, 5298 => 0, 5299 => 0, 5300 => 0, 5301 => 0, 5302 => 1, 5303 => 1, 5304 => 1, 5305 => 1, 5306 => 1, 5307 => 1, 5308 => 1, 5309 => 1, 5310 => 1, 5311 => 1, 5312 => 1, 5313 => 0, 5314 => 0, 5315 => 0, 5316 => 0, 5317 => 0, 5318 => 0, 5319 => 0, 5320 => 0, 5321 => 0, 5322 => 0, 5323 => 0, 5324 => 0, 5325 => 0, 5326 => 0, 5327 => 0, 5328 => 0, 5329 => 0, 5330 => 0, 
5331 => 0, 5332 => 0, 5333 => 0, 5334 => 1, 5335 => 1, 5336 => 1, 5337 => 1, 5338 => 1, 5339 => 1, 5340 => 1, 5341 => 1, 5342 => 1, 5343 => 1, 5344 => 
1, 5345 => 0, 5346 => 0, 5347 => 1, 5348 => 1, 5349 => 1, 5350 => 1, 5351 => 1, 5352 => 1, 5353 => 1, 5354 => 1, 5355 => 1, 5356 => 1, 5357 => 1, 5358 
=> 1, 5359 => 1, 5360 => 1, 5361 => 1, 5362 => 1, 5363 => 1, 5364 => 1, 5365 => 1, 5366 => 1, 5367 => 1, 5368 => 1, 5369 => 1, 5370 => 1, 5371 => 1, 5372 => 1, 5373 => 1, 5374 => 1, 5375 => 1, 5376 => 1, 5377 => 1, 5378 => 1, 5379 => 1, 5380 => 1, 5381 => 1, 5382 => 1, 5383 => 0, 5384 => 0, 5385 => 0, 5386 => 0, 5387 => 0, 5388 => 0, 5389 => 0, 5390 => 0, 5391 => 0, 5392 => 0, 5393 => 0, 5394 => 0, 5395 => 0, 5396 => 0, 5397 => 0, 5398 => 1, 5399 => 1, 5400 => 1, 5401 => 1, 5402 => 1, 5403 => 1, 5404 => 1, 5405 => 1, 5406 => 1, 5407 => 1, 5408 => 1, 5409 => 0, 5410 => 0, 5411 => 0, 5412 => 0, 5413 => 0, 5414 => 0, 5415 => 0, 5416 => 0, 5417 => 0, 5418 => 0, 5419 => 0, 5420 => 0, 5421 => 0, 5422 => 0, 5423 => 0, 5424 => 0, 5425 => 0, 5426 => 0, 5427 => 0, 5428 => 0, 5429 => 0, 5430 => 1, 5431 => 1, 5432 => 1, 5433 => 1, 5434 => 1, 5435 => 1, 5436 => 1, 5437 => 1, 5438 => 1, 5439 => 1, 5440 => 1, 5441 => 0, 5442 => 0, 5443 => 0, 5444 => 0, 5445 => 0, 5446 => 0, 5447 => 0, 5448 => 0, 5449 => 1, 5450 => 1, 5451 => 1, 5452 => 1, 5453 => 1, 5454 => 1, 5455 => 1, 5456 => 1, 5457 => 1, 5458 => 1, 5459 => 1, 5460 => 0, 5461 => 0, 5462 => 0, 5463 => 0, 5464 => 0, 5465 => 0, 5466 => 0, 5467 => 0, 5468 => 0, 5469 => 0, 5470 => 0, 5471 => 0, 5472 => 0, 5473 => 0, 5474 => 1, 5475 => 1, 5476 => 1, 5477 => 1, 5478 => 1, 5479 => 1, 5480 => 1, 5481 => 1, 
5482 => 1, 5483 => 1, 5484 => 1, 5485 => 1, 5486 => 1, 5487 => 1, 5488 => 1, 5489 => 1, 5490 => 1, 5491 => 1, 5492 => 0, 5493 => 0, 5494 => 0, 5495 => 
0, 5496 => 0, 5497 => 0, 5498 => 0, 5499 => 0, 5500 => 1, 5501 => 1, 5502 => 1, 5503 => 1, 5504 => 1, 5505 => 1, 5506 => 1, 5507 => 1, 5508 => 1, 5509 
=> 1, 5510 => 1, 5511 => 0, 5512 => 0, 5513 => 0, 5514 => 0, 5515 => 0, 5516 => 0, 5517 => 0, 5518 => 0, 5519 => 0, 5520 => 0, 5521 => 0, 5522 => 0, 5523 => 0, 5524 => 0, 5525 => 0, 5526 => 0, 5527 => 0, 5528 => 0, 5529 => 0, 5530 => 0, 5531 => 0, 5532 => 1, 5533 => 1, 5534 => 1, 5535 => 1, 5536 => 1, 5537 => 1, 5538 => 1, 5539 => 1, 5540 => 1, 5541 => 1, 5542 => 1, 5543 => 0, 5544 => 0, 5545 => 1, 5546 => 1, 5547 => 1, 5548 => 1, 5549 => 1, 5550 => 1, 5551 => 1, 5552 => 1, 5553 => 1, 5554 => 1, 5555 => 1, 5556 => 1, 5557 => 1, 5558 => 1, 5559 => 1, 5560 => 1, 5561 => 1, 5562 => 1, 5563 => 1, 5564 => 1, 5565 => 1, 5566 => 1, 5567 => 1, 5568 => 1, 5569 => 1, 5570 => 1, 5571 => 1, 5572 => 1, 5573 => 1, 5574 => 1, 5575 => 1, 5576 => 1, 5577 => 1, 5578 => 1, 5579 => 1, 5580 => 1, 5581 => 0, 5582 => 0, 5583 => 0, 5584 => 0, 5585 => 0, 5586 => 0, 5587 => 0, 5588 => 0, 5589 => 0, 5590 => 0, 5591 => 0, 5592 => 0, 5593 => 0, 5594 => 0, 5595 => 0, 5596 => 1, 5597 => 1, 5598 => 1, 5599 => 1, 5600 => 1, 5601 => 1, 5602 => 1, 5603 => 1, 5604 => 1, 5605 => 1, 5606 => 1, 5607 => 0, 5608 => 0, 5609 => 0, 5610 => 0, 5611 => 0, 5612 => 0, 5613 => 0, 5614 => 0, 5615 => 0, 5616 => 0, 5617 => 0, 5618 => 0, 5619 => 0, 5620 => 0, 5621 => 0, 5622 => 0, 5623 => 0, 5624 => 0, 5625 => 0, 5626 => 0, 5627 => 0, 5628 => 1, 5629 => 1, 5630 => 1, 5631 => 1, 5632 => 1, 
5633 => 1, 5634 => 1, 5635 => 1, 5636 => 1, 5637 => 1, 5638 => 1, 5639 => 0, 5640 => 0, 5641 => 0, 5642 => 0, 5643 => 0, 5644 => 0, 5645 => 0, 5646 => 
0, 5647 => 1, 5648 => 1, 5649 => 1, 5650 => 1, 5651 => 1, 5652 => 1, 5653 => 1, 5654 => 1, 5655 => 1, 5656 => 1, 5657 => 1, 5658 => 0, 5659 => 0, 5660 
=> 0, 5661 => 0, 5662 => 0, 5663 => 0, 5664 => 0, 5665 => 0, 5666 => 0, 5667 => 0, 5668 => 0, 5669 => 0, 5670 => 0, 5671 => 0, 5672 => 1, 5673 => 1, 5674 => 1, 5675 => 1, 5676 => 1, 5677 => 1, 5678 => 1, 5679 => 1, 5680 => 1, 5681 => 1, 5682 => 1, 5683 => 1, 5684 => 1, 5685 => 1, 5686 => 1, 5687 => 1, 5688 => 1, 5689 => 1, 5690 => 0, 5691 => 0, 5692 => 0, 5693 => 0, 5694 => 0, 5695 => 0, 5696 => 0, 5697 => 0, 5698 => 1, 5699 => 1, 5700 => 1, 5701 => 1, 5702 => 1, 5703 => 1, 5704 => 1, 5705 => 1, 5706 => 1, 5707 => 1, 5708 => 1, 5709 => 0, 5710 => 0, 5711 => 0, 5712 => 0, 5713 => 0, 5714 => 0, 5715 => 0, 5716 => 0, 5717 => 0, 5718 => 0, 5719 => 0, 5720 => 0, 5721 => 0, 5722 => 0, 5723 => 0, 5724 => 0, 5725 => 0, 5726 => 0, 5727 => 0, 5728 => 0, 5729 => 0, 5730 => 1, 5731 => 1, 5732 => 1, 5733 => 1, 5734 => 1, 5735 => 1, 5736 => 1, 5737 => 1, 5738 => 1, 5739 => 1, 5740 => 1, 5741 => 0, 5742 => 0, 5743 => 1, 5744 => 1, 5745 => 1, 5746 => 1, 5747 => 1, 5748 => 1, 5749 => 1, 5750 => 1, 5751 => 1, 5752 => 1, 5753 => 1, 5754 => 1, 5755 => 1, 5756 => 1, 5757 => 1, 5758 => 1, 5759 => 1, 5760 => 1, 5761 => 1, 5762 => 1, 5763 => 1, 5764 => 1, 5765 => 1, 5766 => 1, 5767 => 1, 5768 => 1, 5769 => 1, 5770 => 1, 5771 => 1, 5772 => 1, 5773 => 1, 5774 => 1, 5775 => 1, 5776 => 1, 5777 => 1, 5778 => 1, 5779 => 0, 5780 => 0, 5781 => 0, 5782 => 0, 5783 => 0, 
5784 => 0, 5785 => 0, 5786 => 0, 5787 => 0, 5788 => 0, 5789 => 0, 5790 => 0, 5791 => 0, 5792 => 0, 5793 => 0, 5794 => 1, 5795 => 1, 5796 => 1, 5797 => 
1, 5798 => 1, 5799 => 1, 5800 => 1, 5801 => 1, 5802 => 1, 5803 => 1, 5804 => 1, 5805 => 0, 5806 => 0, 5807 => 0, 5808 => 0, 5809 => 0, 5810 => 0, 5811 
=> 0, 5812 => 0, 5813 => 0, 5814 => 0, 5815 => 0, 5816 => 0, 5817 => 0, 5818 => 0, 5819 => 0, 5820 => 0, 5821 => 0, 5822 => 0, 5823 => 0, 5824 => 0, 5825 => 0, 5826 => 1, 5827 => 1, 5828 => 1, 5829 => 1, 5830 => 1, 5831 => 1, 5832 => 1, 5833 => 1, 5834 => 1, 5835 => 1, 5836 => 1, 5837 => 0, 5838 => 0, 5839 => 0, 5840 => 0, 5841 => 0, 5842 => 0, 5843 => 0, 5844 => 0, 5845 => 1, 5846 => 1, 5847 => 1, 5848 => 1, 5849 => 1, 5850 => 1, 5851 => 1, 5852 => 1, 5853 => 1, 5854 => 1, 5855 => 1, 5856 => 0, 5857 => 0, 5858 => 0, 5859 => 0, 5860 => 0, 5861 => 0, 5862 => 0, 5863 => 0, 5864 => 0, 5865 => 0, 5866 => 0, 5867 => 0, 5868 => 0, 5869 => 0, 5870 => 1, 5871 => 1, 5872 => 1, 5873 => 1, 5874 => 1, 5875 => 1, 5876 => 1, 5877 => 1, 5878 => 1, 5879 => 1, 5880 => 1, 5881 => 1, 5882 => 1, 5883 => 1, 5884 => 1, 5885 => 1, 5886 => 1, 5887 => 1, 5888 => 0, 5889 => 0, 5890 => 0, 5891 => 0, 5892 => 0, 5893 => 0, 5894 => 0, 5895 => 0, 5896 => 1, 5897 => 1, 5898 => 1, 5899 => 1, 5900 => 1, 5901 => 1, 5902 => 1, 5903 => 1, 5904 => 1, 5905 => 1, 5906 => 1, 5907 => 0, 5908 => 0, 5909 => 0, 5910 => 0, 5911 => 0, 5912 => 0, 5913 => 0, 5914 => 0, 5915 => 0, 5916 => 0, 5917 => 0, 5918 => 0, 5919 => 0, 5920 => 0, 5921 => 0, 5922 => 0, 5923 => 0, 5924 => 0, 5925 => 0, 5926 => 0, 5927 => 0, 5928 => 1, 5929 => 1, 5930 => 1, 5931 => 1, 5932 => 1, 5933 => 1, 5934 => 1, 
5935 => 1, 5936 => 1, 5937 => 1, 5938 => 1, 5939 => 0, 5940 => 0, 5941 => 1, 5942 => 1, 5943 => 1, 5944 => 1, 5945 => 1, 5946 => 1, 5947 => 1, 5948 => 
1, 5949 => 1, 5950 => 1, 5951 => 1, 5952 => 1, 5953 => 1, 5954 => 1, 5955 => 1, 5956 => 1, 5957 => 1, 5958 => 1, 5959 => 1, 5960 => 1, 5961 => 1, 5962 
=> 1, 5963 => 1, 5964 => 1, 5965 => 1, 5966 => 1, 5967 => 1, 5968 => 1, 5969 => 1, 5970 => 1, 5971 => 1, 5972 => 1, 5973 => 1, 5974 => 1, 5975 => 1, 5976 => 1, 5977 => 0, 5978 => 0, 5979 => 0, 5980 => 0, 5981 => 0, 5982 => 0, 5983 => 0, 5984 => 0, 5985 => 0, 5986 => 0, 5987 => 0, 5988 => 0, 5989 => 0, 5990 => 0, 5991 => 0, 5992 => 1, 5993 => 1, 5994 => 1, 5995 => 1, 5996 => 1, 5997 => 1, 5998 => 1, 5999 => 1, 6000 => 1, 6001 => 1, 6002 => 1, 6003 => 0, 6004 => 0, 6005 => 0, 6006 => 0, 6007 => 0, 6008 => 0, 6009 => 0, 6010 => 0, 6011 => 0, 6012 => 0, 6013 => 0, 6014 => 0, 6015 => 0, 6016 => 0, 6017 => 0, 6018 => 0, 6019 => 0, 6020 => 0, 6021 => 0, 6022 => 0, 6023 => 0, 6024 => 1, 6025 => 1, 6026 => 1, 6027 => 1, 6028 => 1, 6029 => 1, 6030 => 1, 6031 => 1, 6032 => 1, 6033 => 1, 6034 => 1, 6035 => 0, 6036 => 0, 6037 => 0, 6038 => 0, 6039 => 0, 6040 => 0, 6041 => 0, 6042 => 0, 6043 => 1, 6044 => 1, 6045 => 1, 6046 => 1, 6047 => 1, 6048 => 1, 6049 => 1, 6050 => 1, 6051 => 1, 6052 => 1, 6053 => 1, 6054 => 0, 6055 => 0, 6056 => 0, 6057 => 0, 6058 => 0, 6059 => 0, 6060 => 0, 6061 => 0, 6062 => 0, 6063 => 0, 6064 => 0, 6065 => 0, 6066 => 0, 6067 => 0, 6068 => 1, 6069 => 1, 6070 => 1, 6071 => 1, 6072 => 1, 6073 => 1, 6074 => 1, 6075 => 1, 6076 => 1, 6077 => 1, 6078 => 1, 6079 => 1, 6080 => 1, 6081 => 1, 6082 => 1, 6083 => 1, 6084 => 1, 6085 => 1, 
6086 => 0, 6087 => 0, 6088 => 0, 6089 => 0, 6090 => 0, 6091 => 0, 6092 => 0, 6093 => 0, 6094 => 1, 6095 => 1, 6096 => 1, 6097 => 1, 6098 => 1, 6099 => 
1, 6100 => 1, 6101 => 1, 6102 => 1, 6103 => 1, 6104 => 1, 6105 => 0, 6106 => 0, 6107 => 0, 6108 => 0, 6109 => 0, 6110 => 0, 6111 => 0, 6112 => 0, 6113 
=> 0, 6114 => 0, 6115 => 0, 6116 => 0, 6117 => 0, 6118 => 0, 6119 => 0, 6120 => 0, 6121 => 0, 6122 => 0, 6123 => 0, 6124 => 0, 6125 => 0, 6126 => 1, 6127 => 1, 6128 => 1, 6129 => 1, 6130 => 1, 6131 => 1, 6132 => 1, 6133 => 1, 6134 => 1, 6135 => 1, 6136 => 1, 6137 => 0, 6138 => 0, 6139 => 1, 6140 => 1, 6141 => 1, 6142 => 1, 6143 => 1, 6144 => 1, 6145 => 1, 6146 => 1, 6147 => 1, 6148 => 1, 6149 => 1, 6150 => 1, 6151 => 0, 6152 => 0, 6153 => 0, 6154 => 0, 6155 => 0, 6156 => 0, 6157 => 0, 6158 => 0, 6159 => 0, 6160 => 0, 6161 => 0, 6162 => 0, 6163 => 0, 6164 => 0, 6165 => 0, 6166 => 0, 6167 => 0, 6168 => 0, 6169 => 0, 6170 => 0, 6171 => 0, 6172 => 0, 6173 => 0, 6174 => 0, 6175 => 0, 6176 => 0, 6177 => 0, 6178 => 0, 6179 => 0, 6180 => 0, 6181 => 0, 6182 => 0, 6183 => 0, 6184 => 0, 6185 => 0, 6186 => 0, 6187 => 0, 6188 => 0, 6189 => 0, 6190 => 1, 6191 => 1, 6192 => 1, 6193 => 1, 6194 => 1, 6195 => 1, 6196 => 1, 6197 => 1, 6198 => 1, 6199 => 1, 6200 => 1, 6201 => 0, 6202 => 0, 6203 => 0, 6204 => 0, 6205 => 0, 6206 => 0, 6207 => 0, 6208 => 0, 6209 => 0, 6210 => 0, 6211 => 0, 6212 => 0, 6213 => 0, 6214 => 0, 6215 => 0, 6216 => 0, 6217 => 0, 6218 => 0, 6219 => 0, 6220 => 0, 6221 => 0, 6222 => 1, 6223 => 1, 6224 => 1, 6225 => 1, 6226 => 1, 6227 => 1, 6228 => 1, 6229 => 1, 6230 => 1, 6231 => 1, 6232 => 1, 6233 => 0, 6234 => 0, 6235 => 0, 6236 => 0, 
6237 => 0, 6238 => 0, 6239 => 0, 6240 => 0, 6241 => 1, 6242 => 1, 6243 => 1, 6244 => 1, 6245 => 1, 6246 => 1, 6247 => 1, 6248 => 1, 6249 => 1, 6250 => 
1, 6251 => 1, 6252 => 0, 6253 => 0, 6254 => 0, 6255 => 0, 6256 => 0, 6257 => 0, 6258 => 0, 6259 => 0, 6260 => 0, 6261 => 0, 6262 => 0, 6263 => 0, 6264 
=> 0, 6265 => 0, 6266 => 1, 6267 => 0, 6268 => 0, 6269 => 0, 6270 => 0, 6271 => 0, 6272 => 1, 6273 => 1, 6274 => 1, 6275 => 1, 6276 => 1, 6277 => 1, 6278 => 1, 6279 => 1, 6280 => 1, 6281 => 1, 6282 => 1, 6283 => 1, 6284 => 0, 6285 => 0, 6286 => 0, 6287 => 0, 6288 => 0, 6289 => 0, 6290 => 0, 6291 => 0, 6292 => 1, 6293 => 1, 6294 => 1, 6295 => 1, 6296 => 1, 6297 => 1, 6298 => 1, 6299 => 1, 6300 => 1, 6301 => 1, 6302 => 1, 6303 => 0, 6304 => 0, 6305 => 0, 6306 => 0, 6307 => 0, 6308 => 0, 6309 => 0, 6310 => 0, 6311 => 0, 6312 => 0, 6313 => 0, 6314 => 0, 6315 => 0, 6316 => 0, 6317 => 0, 6318 => 0, 6319 => 0, 6320 => 0, 6321 => 0, 6322 => 0, 6323 => 0, 6324 => 1, 6325 => 1, 6326 => 1, 6327 => 1, 6328 => 1, 6329 => 1, 6330 => 1, 6331 => 1, 6332 => 1, 6333 => 1, 6334 => 1, 6335 => 0, 6336 => 0, 6337 => 1, 6338 => 1, 6339 => 1, 6340 => 1, 6341 => 1, 6342 => 1, 6343 => 1, 6344 => 1, 6345 => 1, 6346 => 1, 6347 => 1, 6348 => 0, 6349 => 0, 6350 => 0, 6351 => 0, 6352 => 0, 6353 => 0, 6354 => 0, 6355 => 0, 6356 => 0, 6357 => 0, 6358 => 0, 6359 => 0, 6360 => 0, 6361 => 0, 6362 => 0, 6363 => 0, 6364 => 0, 6365 => 0, 6366 => 0, 6367 => 0, 6368 => 0, 6369 => 0, 6370 => 0, 6371 => 0, 6372 => 0, 6373 => 0, 6374 => 0, 6375 => 0, 6376 => 0, 6377 => 0, 6378 => 0, 6379 => 0, 6380 => 0, 6381 => 0, 6382 => 0, 6383 => 0, 6384 => 0, 6385 => 0, 6386 => 0, 6387 => 0, 
6388 => 1, 6389 => 1, 6390 => 1, 6391 => 1, 6392 => 1, 6393 => 1, 6394 => 1, 6395 => 1, 6396 => 1, 6397 => 1, 6398 => 1, 6399 => 0, 6400 => 0, 6401 => 
0, 6402 => 0, 6403 => 0, 6404 => 0, 6405 => 0, 6406 => 0, 6407 => 0, 6408 => 0, 6409 => 0, 6410 => 0, 6411 => 0, 6412 => 0, 6413 => 0, 6414 => 0, 6415 
=> 0, 6416 => 0, 6417 => 0, 6418 => 0, 6419 => 0, 6420 => 1, 6421 => 1, 6422 => 1, 6423 => 1, 6424 => 1, 6425 => 1, 6426 => 1, 6427 => 1, 6428 => 1, 6429 => 1, 6430 => 1, 6431 => 0, 6432 => 0, 6433 => 0, 6434 => 0, 6435 => 0, 6436 => 0, 6437 => 0, 6438 => 0, 6439 => 1, 6440 => 1, 6441 => 1, 6442 => 1, 6443 => 1, 6444 => 1, 6445 => 1, 6446 => 1, 6447 => 1, 6448 => 1, 6449 => 1, 6450 => 0, 6451 => 0, 6452 => 0, 6453 => 0, 6454 => 0, 6455 => 0, 6456 => 0, 6457 => 0, 6458 => 0, 6459 => 0, 6460 => 0, 6461 => 0, 6462 => 0, 6463 => 0, 6464 => 0, 6465 => 0, 6466 => 0, 6467 => 0, 6468 => 0, 6469 => 0, 6470 => 0, 6471 => 1, 6472 => 1, 6473 => 1, 6474 => 1, 6475 => 1, 6476 => 1, 6477 => 1, 6478 => 1, 6479 => 1, 6480 => 1, 6481 => 1, 6482 => 0, 6483 => 0, 6484 => 0, 6485 => 0, 6486 => 0, 6487 => 0, 6488 => 0, 6489 => 0, 6490 => 1, 6491 => 1, 6492 => 1, 6493 => 1, 6494 => 1, 6495 => 1, 6496 => 1, 6497 => 1, 6498 => 1, 6499 => 1, 6500 => 1, 6501 => 0, 6502 => 0, 6503 => 0, 6504 => 0, 6505 => 0, 6506 => 0, 6507 => 0, 6508 => 0, 6509 => 0, 6510 => 0, 6511 => 0, 6512 => 0, 6513 => 0, 6514 => 0, 6515 => 0, 6516 => 0, 6517 => 0, 6518 => 0, 6519 => 0, 6520 => 0, 6521 => 0, 6522 => 1, 6523 => 1, 6524 => 1, 6525 => 1, 6526 => 1, 6527 => 1, 6528 => 1, 6529 => 1, 6530 => 1, 6531 => 1, 6532 => 1, 6533 => 0, 6534 => 0, 6535 => 1, 6536 => 1, 6537 => 1, 6538 => 1, 
6539 => 1, 6540 => 1, 6541 => 1, 6542 => 1, 6543 => 1, 6544 => 1, 6545 => 1, 6546 => 0, 6547 => 0, 6548 => 0, 6549 => 0, 6550 => 0, 6551 => 0, 6552 => 
0, 6553 => 0, 6554 => 0, 6555 => 0, 6556 => 0, 6557 => 0, 6558 => 0, 6559 => 0, 6560 => 0, 6561 => 0, 6562 => 0, 6563 => 0, 6564 => 0, 6565 => 0, 6566 
=> 0, 6567 => 0, 6568 => 0, 6569 => 0, 6570 => 0, 6571 => 0, 6572 => 0, 6573 => 0, 6574 => 0, 6575 => 0, 6576 => 0, 6577 => 0, 6578 => 0, 6579 => 0, 6580 => 0, 6581 => 0, 6582 => 0, 6583 => 0, 6584 => 0, 6585 => 0, 6586 => 1, 6587 => 1, 6588 => 1, 6589 => 1, 6590 => 1, 6591 => 1, 6592 => 1, 6593 => 1, 6594 => 1, 6595 => 1, 6596 => 1, 6597 => 0, 6598 => 0, 6599 => 0, 6600 => 0, 6601 => 0, 6602 => 0, 6603 => 0, 6604 => 0, 6605 => 0, 6606 => 0, 6607 => 0, 6608 => 0, 6609 => 0, 6610 => 0, 6611 => 0, 6612 => 0, 6613 => 0, 6614 => 0, 6615 => 0, 6616 => 0, 6617 => 0, 6618 => 1, 6619 => 1, 6620 => 1, 6621 => 1, 6622 => 1, 6623 => 1, 6624 => 1, 6625 => 1, 6626 => 1, 6627 => 1, 6628 => 1, 6629 => 0, 6630 => 0, 6631 => 0, 6632 => 0, 6633 => 0, 6634 => 0, 6635 => 0, 6636 => 0, 6637 => 1, 6638 => 1, 6639 => 1, 6640 => 1, 6641 => 1, 6642 => 1, 6643 => 1, 6644 => 1, 6645 => 1, 6646 => 1, 6647 => 1, 6648 => 0, 6649 => 0, 6650 => 0, 6651 => 0, 6652 => 0, 6653 => 0, 6654 => 0, 6655 => 0, 6656 => 0, 6657 => 0, 6658 => 0, 6659 => 0, 6660 => 0, 6661 => 0, 6662 => 0, 6663 => 0, 6664 => 0, 6665 => 0, 6666 => 0, 6667 => 0, 6668 => 0, 6669 => 1, 6670 => 1, 6671 => 1, 6672 => 1, 6673 => 1, 6674 => 1, 6675 => 1, 6676 => 1, 6677 => 1, 6678 => 1, 6679 => 1, 6680 => 0, 6681 => 0, 6682 => 0, 6683 => 0, 6684 => 0, 6685 => 0, 6686 => 0, 6687 => 0, 6688 => 1, 6689 => 1, 
6690 => 1, 6691 => 1, 6692 => 1, 6693 => 1, 6694 => 1, 6695 => 1, 6696 => 1, 6697 => 1, 6698 => 1, 6699 => 0, 6700 => 0, 6701 => 0, 6702 => 0, 6703 => 
0, 6704 => 0, 6705 => 0, 6706 => 0, 6707 => 0, 6708 => 0, 6709 => 0, 6710 => 0, 6711 => 0, 6712 => 0, 6713 => 0, 6714 => 0, 6715 => 0, 6716 => 0, 6717 
=> 0, 6718 => 0, 6719 => 0, 6720 => 1, 6721 => 1, 6722 => 1, 6723 => 1, 6724 => 1, 6725 => 1, 6726 => 1, 6727 => 1, 6728 => 1, 6729 => 1, 6730 => 1, 6731 => 0, 6732 => 0, 6733 => 1, 6734 => 1, 6735 => 1, 6736 => 1, 6737 => 1, 6738 => 1, 6739 => 1, 6740 => 1, 6741 => 1, 6742 => 1, 6743 => 1, 6744 => 0, 6745 => 0, 6746 => 0, 6747 => 0, 6748 => 0, 6749 => 0, 6750 => 0, 6751 => 0, 6752 => 0, 6753 => 0, 6754 => 0, 6755 => 0, 6756 => 0, 6757 => 0, 6758 => 0, 6759 => 0, 6760 => 0, 6761 => 0, 6762 => 0, 6763 => 0, 6764 => 0, 6765 => 0, 6766 => 0, 6767 => 0, 6768 => 0, 6769 => 0, 6770 => 0, 6771 => 0, 6772 => 0, 6773 => 0, 6774 => 0, 6775 => 0, 6776 => 0, 6777 => 0, 6778 => 0, 6779 => 0, 6780 => 0, 6781 => 0, 6782 => 0, 6783 => 0, 6784 => 1, 6785 => 1, 6786 => 1, 6787 => 1, 6788 => 1, 6789 => 1, 6790 => 1, 6791 => 1, 6792 => 1, 6793 => 1, 6794 => 1, 6795 => 0, 6796 => 0, 6797 => 0, 6798 => 0, 6799 => 0, 6800 => 0, 6801 => 0, 6802 => 0, 6803 => 0, 6804 => 0, 6805 => 0, 6806 => 0, 6807 => 0, 6808 => 0, 6809 => 0, 6810 => 0, 6811 => 0, 6812 => 0, 6813 => 0, 6814 => 0, 6815 => 0, 6816 => 1, 6817 => 1, 6818 => 1, 6819 => 1, 6820 => 1, 6821 => 1, 6822 => 1, 6823 => 1, 6824 => 1, 6825 => 1, 6826 => 1, 6827 => 0, 6828 => 0, 6829 => 0, 6830 => 0, 6831 => 0, 6832 => 0, 6833 => 0, 6834 => 0, 6835 => 1, 6836 => 1, 6837 => 1, 6838 => 1, 6839 => 1, 6840 => 1, 
6841 => 1, 6842 => 1, 6843 => 1, 6844 => 1, 6845 => 1, 6846 => 0, 6847 => 0, 6848 => 0, 6849 => 0, 6850 => 0, 6851 => 0, 6852 => 0, 6853 => 0, 6854 => 
0, 6855 => 0, 6856 => 0, 6857 => 0, 6858 => 0, 6859 => 0, 6860 => 0, 6861 => 0, 6862 => 0, 6863 => 0, 6864 => 0, 6865 => 0, 6866 => 0, 6867 => 1, 6868 
=> 1, 6869 => 1, 6870 => 1, 6871 => 1, 6872 => 1, 6873 => 1, 6874 => 1, 6875 => 1, 6876 => 1, 6877 => 1, 6878 => 0, 6879 => 0, 6880 => 0, 6881 => 0, 6882 => 0, 6883 => 0, 6884 => 0, 6885 => 0, 6886 => 1, 6887 => 1, 6888 => 1, 6889 => 1, 6890 => 1, 6891 => 1, 6892 => 1, 6893 => 1, 6894 => 1, 6895 => 1, 6896 => 1, 6897 => 0, 6898 => 0, 6899 => 0, 6900 => 0, 6901 => 0, 6902 => 0, 6903 => 0, 6904 => 0, 6905 => 0, 6906 => 0, 6907 => 0, 6908 => 0, 6909 => 0, 6910 => 0, 6911 => 0, 6912 => 0, 6913 => 0, 6914 => 0, 6915 => 0, 6916 => 0, 6917 => 0, 6918 => 1, 6919 => 1, 6920 => 1, 6921 => 1, 6922 => 1, 6923 => 1, 6924 => 1, 6925 => 1, 6926 => 1, 6927 => 1, 6928 => 1, 6929 => 0, 6930 => 0, 6931 => 1, 6932 => 1, 6933 => 1, 6934 => 1, 6935 => 1, 6936 => 1, 6937 => 1, 6938 => 1, 6939 => 1, 6940 => 1, 6941 => 1, 6942 => 0, 6943 => 0, 6944 => 0, 6945 => 0, 6946 => 0, 6947 => 0, 6948 => 0, 6949 => 0, 6950 => 0, 6951 => 0, 6952 => 0, 6953 => 0, 6954 => 0, 6955 => 0, 6956 => 0, 6957 => 0, 6958 => 0, 6959 => 0, 6960 => 0, 6961 => 0, 6962 => 0, 6963 => 0, 6964 => 0, 6965 => 0, 6966 => 0, 6967 => 0, 6968 => 0, 6969 => 0, 6970 => 0, 6971 => 0, 6972 => 0, 6973 => 0, 6974 => 0, 6975 => 0, 6976 => 0, 6977 => 0, 6978 => 0, 6979 => 0, 6980 => 0, 6981 => 0, 6982 => 1, 6983 => 1, 6984 => 1, 6985 => 1, 6986 => 1, 6987 => 1, 6988 => 1, 6989 => 1, 6990 => 1, 6991 => 1, 
6992 => 1, 6993 => 0, 6994 => 0, 6995 => 0, 6996 => 0, 6997 => 0, 6998 => 0, 6999 => 0, 7000 => 0, 7001 => 0, 7002 => 0, 7003 => 0, 7004 => 0, 7005 => 
0, 7006 => 0, 7007 => 0, 7008 => 0, 7009 => 0, 7010 => 0, 7011 => 0, 7012 => 0, 7013 => 0, 7014 => 1, 7015 => 1, 7016 => 1, 7017 => 1, 7018 => 1, 7019 
=> 1, 7020 => 1, 7021 => 1, 7022 => 1, 7023 => 1, 7024 => 1, 7025 => 0, 7026 => 0, 7027 => 0, 7028 => 0, 7029 => 0, 7030 => 0, 7031 => 0, 7032 => 0, 7033 => 1, 7034 => 1, 7035 => 1, 7036 => 1, 7037 => 1, 7038 => 1, 7039 => 1, 7040 => 1, 7041 => 1, 7042 => 1, 7043 => 1, 7044 => 0, 7045 => 0, 7046 => 0, 7047 => 0, 7048 => 0, 7049 => 0, 7050 => 0, 7051 => 0, 7052 => 0, 7053 => 0, 7054 => 0, 7055 => 0, 7056 => 0, 7057 => 0, 7058 => 0, 7059 => 0, 7060 => 0, 7061 => 0, 7062 => 0, 7063 => 0, 7064 => 0, 7065 => 1, 7066 => 1, 7067 => 1, 7068 => 1, 7069 => 1, 7070 => 1, 7071 => 1, 7072 => 1, 7073 => 1, 7074 => 1, 7075 => 1, 7076 => 0, 7077 => 0, 7078 => 0, 7079 => 0, 7080 => 0, 7081 => 0, 7082 => 0, 7083 => 0, 7084 => 1, 7085 => 1, 7086 => 1, 7087 => 1, 7088 => 1, 7089 => 1, 7090 => 1, 7091 => 1, 7092 => 1, 7093 => 1, 7094 => 1, 7095 => 0, 7096 => 0, 7097 => 0, 7098 => 0, 7099 => 0, 7100 => 0, 7101 => 0, 7102 => 0, 7103 => 0, 7104 => 0, 7105 => 0, 7106 => 0, 7107 => 0, 7108 => 0, 7109 => 0, 7110 => 0, 7111 => 0, 7112 => 0, 7113 => 0, 7114 => 0, 7115 => 0, 7116 => 1, 7117 => 1, 7118 => 1, 7119 => 1, 7120 => 1, 7121 => 1, 7122 => 1, 7123 => 1, 7124 => 1, 7125 => 1, 7126 => 1, 7127 => 0, 7128 => 0, 7129 => 1, 7130 => 1, 7131 => 1, 7132 => 1, 7133 => 1, 7134 => 1, 7135 => 1, 7136 => 1, 7137 => 1, 7138 => 1, 7139 => 1, 7140 => 0, 7141 => 0, 7142 => 0, 
7143 => 0, 7144 => 0, 7145 => 0, 7146 => 0, 7147 => 0, 7148 => 0, 7149 => 0, 7150 => 0, 7151 => 0, 7152 => 0, 7153 => 0, 7154 => 0, 7155 => 0, 7156 => 
0, 7157 => 0, 7158 => 0, 7159 => 0, 7160 => 0, 7161 => 0, 7162 => 0, 7163 => 0, 7164 => 0, 7165 => 0, 7166 => 0, 7167 => 0, 7168 => 0, 7169 => 0, 7170 
=> 0, 7171 => 0, 7172 => 0, 7173 => 0, 7174 => 0, 7175 => 0, 7176 => 0, 7177 => 0, 7178 => 0, 7179 => 0, 7180 => 1, 7181 => 1, 7182 => 1, 7183 => 1, 7184 => 1, 7185 => 1, 7186 => 1, 7187 => 1, 7188 => 1, 7189 => 1, 7190 => 1, 7191 => 0, 7192 => 0, 7193 => 0, 7194 => 0, 7195 => 0, 7196 => 0, 7197 => 0, 7198 => 0, 7199 => 0, 7200 => 0, 7201 => 0, 7202 => 0, 7203 => 0, 7204 => 0, 7205 => 0, 7206 => 0, 7207 => 0, 7208 => 0, 7209 => 0, 7210 => 0, 7211 => 0, 7212 => 1, 7213 => 1, 7214 => 1, 7215 => 1, 7216 => 1, 7217 => 1, 7218 => 1, 7219 => 1, 7220 => 1, 7221 => 1, 7222 => 1, 7223 => 0, 7224 => 0, 7225 => 0, 7226 => 0, 7227 => 0, 7228 => 0, 7229 => 0, 7230 => 0, 7231 => 1, 7232 => 1, 7233 => 1, 7234 => 1, 7235 => 1, 7236 => 1, 7237 => 1, 7238 => 1, 7239 => 1, 7240 => 1, 7241 => 1, 7242 => 0, 7243 => 0, 7244 => 0, 7245 => 0, 7246 => 0, 7247 => 0, 7248 => 0, 7249 => 0, 7250 => 0, 7251 => 0, 7252 => 0, 7253 => 0, 7254 => 0, 7255 => 0, 7256 => 0, 7257 => 0, 7258 => 0, 7259 => 0, 7260 => 0, 7261 => 0, 7262 => 0, 7263 => 1, 7264 => 1, 7265 => 1, 7266 => 1, 7267 => 1, 7268 => 1, 7269 => 1, 7270 => 1, 7271 => 1, 7272 => 1, 7273 => 1, 7274 => 0, 7275 => 0, 7276 => 0, 7277 => 0, 7278 => 0, 7279 => 0, 7280 => 0, 7281 => 0, 7282 => 1, 7283 => 1, 7284 => 1, 7285 => 1, 7286 => 1, 7287 => 1, 7288 => 1, 7289 => 1, 7290 => 1, 7291 => 1, 7292 => 1, 7293 => 0, 
7294 => 0, 7295 => 0, 7296 => 0, 7297 => 0, 7298 => 0, 7299 => 0, 7300 => 0, 7301 => 0, 7302 => 0, 7303 => 0, 7304 => 0, 7305 => 0, 7306 => 0, 7307 => 
0, 7308 => 0, 7309 => 0, 7310 => 0, 7311 => 0, 7312 => 0, 7313 => 0, 7314 => 1, 7315 => 1, 7316 => 1, 7317 => 1, 7318 => 1, 7319 => 1, 7320 => 1, 7321 
=> 1, 7322 => 1, 7323 => 1, 7324 => 1, 7325 => 0, 7326 => 0, 7327 => 1, 7328 => 1, 7329 => 1, 7330 => 1, 7331 => 1, 7332 => 1, 7333 => 1, 7334 => 1, 7335 => 1, 7336 => 1, 7337 => 1, 7338 => 0, 7339 => 0, 7340 => 0, 7341 => 0, 7342 => 0, 7343 => 0, 7344 => 0, 7345 => 0, 7346 => 0, 7347 => 0, 7348 => 0, 7349 => 0, 7350 => 0, 7351 => 0, 7352 => 0, 7353 => 0, 7354 => 0, 7355 => 0, 7356 => 0, 7357 => 0, 7358 => 0, 7359 => 0, 7360 => 0, 7361 => 0, 7362 => 0, 7363 => 0, 7364 => 0, 7365 => 0, 7366 => 0, 7367 => 0, 7368 => 0, 7369 => 0, 7370 => 0, 7371 => 0, 7372 => 0, 7373 => 0, 7374 => 0, 7375 => 0, 7376 => 0, 7377 => 0, 7378 => 1, 7379 => 1, 7380 => 1, 7381 => 1, 7382 => 1, 7383 => 1, 7384 => 1, 7385 => 1, 7386 => 1, 7387 => 1, 7388 => 1, 7389 => 0, 7390 => 0, 7391 => 0, 7392 => 0, 7393 => 0, 7394 => 0, 7395 => 0, 7396 => 0, 7397 => 0, 7398 => 0, 7399 => 0, 7400 => 0, 7401 => 0, 7402 => 0, 7403 => 0, 7404 => 0, 7405 => 0, 7406 => 0, 7407 => 0, 7408 => 0, 7409 => 0, 7410 => 1, 7411 => 1, 7412 => 1, 7413 => 1, 7414 => 1, 7415 => 1, 7416 => 1, 7417 => 1, 7418 => 1, 7419 => 1, 7420 => 1, 7421 => 0, 7422 => 0, 7423 => 0, 7424 => 0, 7425 => 0, 7426 => 0, 7427 => 0, 7428 => 0, 7429 => 1, 7430 => 1, 7431 => 1, 7432 => 1, 7433 => 1, 7434 => 1, 7435 => 1, 7436 => 1, 7437 => 1, 7438 => 1, 7439 => 1, 7440 => 0, 7441 => 0, 7442 => 0, 7443 => 0, 7444 => 0, 
7445 => 0, 7446 => 0, 7447 => 0, 7448 => 0, 7449 => 0, 7450 => 0, 7451 => 0, 7452 => 0, 7453 => 0, 7454 => 0, 7455 => 0, 7456 => 0, 7457 => 0, 7458 => 
0, 7459 => 0, 7460 => 0, 7461 => 1, 7462 => 1, 7463 => 1, 7464 => 1, 7465 => 1, 7466 => 1, 7467 => 1, 7468 => 1, 7469 => 1, 7470 => 1, 7471 => 1, 7472 
=> 0, 7473 => 0, 7474 => 0, 7475 => 0, 7476 => 0, 7477 => 0, 7478 => 0, 7479 => 0, 7480 => 1, 7481 => 1, 7482 => 1, 7483 => 1, 7484 => 1, 7485 => 1, 7486 => 1, 7487 => 1, 7488 => 1, 7489 => 1, 7490 => 1, 7491 => 0, 7492 => 0, 7493 => 0, 7494 => 0, 7495 => 0, 7496 => 0, 7497 => 0, 7498 => 0, 7499 => 0, 7500 => 0, 7501 => 0, 7502 => 0, 7503 => 0, 7504 => 0, 7505 => 0, 7506 => 0, 7507 => 0, 7508 => 0, 7509 => 0, 7510 => 0, 7511 => 0, 7512 => 1, 7513 => 1, 7514 => 1, 7515 => 1, 7516 => 1, 7517 => 1, 7518 => 1, 7519 => 1, 7520 => 1, 7521 => 1, 7522 => 1, 7523 => 0, 7524 => 0, 7525 => 1, 7526 => 1, 7527 => 1, 7528 => 1, 7529 => 1, 7530 => 1, 7531 => 1, 7532 => 1, 7533 => 1, 7534 => 1, 7535 => 1, 7536 => 0, 7537 => 0, 7538 => 0, 7539 => 0, 7540 => 0, 7541 => 0, 7542 => 0, 7543 => 0, 7544 => 0, 7545 => 0, 7546 => 0, 7547 => 0, 7548 => 0, 7549 => 0, 7550 => 0, 7551 => 0, 7552 => 0, 7553 => 0, 7554 => 0, 7555 => 0, 7556 => 0, 7557 => 0, 7558 => 0, 7559 => 0, 7560 => 0, 7561 => 0, 7562 => 0, 7563 => 0, 7564 => 0, 7565 => 0, 7566 => 0, 7567 => 0, 7568 => 0, 7569 => 0, 7570 => 0, 7571 => 0, 7572 => 0, 7573 => 0, 7574 => 0, 7575 => 0, 7576 => 0, 7577 => 0, 7578 => 0, 7579 => 0, 7580 => 0, 7581 => 0, 7582 => 1, 7583 => 1, 7584 => 1, 7585 => 1, 7586 => 1, 7587 => 0, 7588 => 0, 7589 => 0, 7590 => 0, 7591 => 0, 7592 => 0, 7593 => 0, 7594 => 0, 7595 => 0, 
7596 => 0, 7597 => 0, 7598 => 0, 7599 => 0, 7600 => 0, 7601 => 0, 7602 => 0, 7603 => 0, 7604 => 0, 7605 => 0, 7606 => 0, 7607 => 0, 7608 => 1, 7609 => 
1, 7610 => 1, 7611 => 1, 7612 => 1, 7613 => 0, 7614 => 0, 7615 => 0, 7616 => 0, 7617 => 0, 7618 => 0, 7619 => 0, 7620 => 0, 7621 => 0, 7622 => 0, 7623 
=> 0, 7624 => 0, 7625 => 0, 7626 => 0, 7627 => 1, 7628 => 1, 7629 => 1, 7630 => 1, 7631 => 1, 7632 => 1, 7633 => 1, 7634 => 1, 7635 => 1, 7636 => 1, 7637 => 1, 7638 => 0, 7639 => 0, 7640 => 0, 7641 => 0, 7642 => 0, 7643 => 0, 7644 => 0, 7645 => 0, 7646 => 0, 7647 => 0, 7648 => 0, 7649 => 0, 7650 => 0, 7651 => 0, 7652 => 0, 7653 => 0, 7654 => 0, 7655 => 0, 7656 => 0, 7657 => 0, 7658 => 0, 7659 => 1, 7660 => 1, 7661 => 1, 7662 => 1, 7663 => 1, 7664 => 1, 7665 => 1, 7666 => 1, 7667 => 1, 7668 => 1, 7669 => 1, 7670 => 0, 7671 => 0, 7672 => 0, 7673 => 0, 7674 => 0, 7675 => 0, 7676 => 0, 7677 => 0, 7678 => 0, 7679 => 0, 7680 => 0, 7681 => 0, 7682 => 0, 7683 => 0, 7684 => 1, 7685 => 1, 7686 => 1, 7687 => 1, 7688 => 1, 7689 => 0, 7690 => 0, 7691 => 0, 7692 => 0, 7693 => 0, 7694 => 0, 7695 => 0, 7696 => 0, 7697 => 0, 7698 => 0, 7699 => 0, 7700 => 0, 7701 => 0, 7702 => 0, 7703 => 0, 7704 => 0, 7705 => 0, 7706 => 0, 7707 => 0, 7708 => 0, 7709 => 0, 7710 => 1, 7711 => 1, 7712 => 1, 7713 => 1, 7714 => 1, 7715 => 0, 7716 => 0, 7717 => 0, 7718 => 0, 7719 => 0, 7720 => 0, 7721 => 0, 7722 => 0, 7723 => 1, 7724 => 1, 7725 => 1, 7726 => 1, 7727 => 1, 7728 => 1, 7729 => 1, 7730 => 1, 7731 => 1, 7732 => 1, 7733 => 1, 7734 => 0, 7735 => 0, 7736 => 0, 7737 => 0, 7738 => 0, 7739 => 0, 7740 => 0, 7741 => 0, 7742 => 0, 7743 => 0, 7744 => 0, 7745 => 0, 7746 => 0, 
7747 => 0, 7748 => 0, 7749 => 0, 7750 => 0, 7751 => 0, 7752 => 0, 7753 => 0, 7754 => 0, 7755 => 0, 7756 => 0, 7757 => 0, 7758 => 0, 7759 => 0, 7760 => 
0, 7761 => 0, 7762 => 0, 7763 => 0, 7764 => 0, 7765 => 0, 7766 => 0, 7767 => 0, 7768 => 0, 7769 => 0, 7770 => 0, 7771 => 0, 7772 => 0, 7773 => 0, 7774 
=> 0, 7775 => 0, 7776 => 0, 7777 => 0, 7778 => 0, 7779 => 0, 7780 => 1, 7781 => 1, 7782 => 1, 7783 => 1, 7784 => 1, 7785 => 1, 7786 => 1, 7787 => 1, 7788 => 1, 7789 => 1, 7790 => 1, 7791 => 1, 7792 => 1, 7793 => 1, 7794 => 1, 7795 => 1, 7796 => 1, 7797 => 1, 7798 => 1, 7799 => 1, 7800 => 1, 7801 => 1, 7802 => 1, 7803 => 1, 7804 => 1, 7805 => 1, 7806 => 1, 7807 => 1, 7808 => 1, 7809 => 1, 7810 => 1, 7811 => 0, 7812 => 0, 7813 => 0, 7814 => 0, 7815 => 0, 7816 => 0, 7817 => 0, 7818 => 0, 7819 => 0, 7820 => 0, 7821 => 0, 7822 => 0, 7823 => 0, 7824 => 0, 7825 => 1, 7826 => 1, 7827 => 1, 7828 => 1, 7829 => 1, 7830 => 1, 7831 => 1, 7832 => 1, 7833 => 1, 7834 => 1, 7835 => 1, 7836 => 0, 7837 => 0, 7838 => 0, 7839 => 0, 7840 => 0, 7841 => 0, 7842 => 0, 7843 => 0, 7844 => 0, 7845 => 0, 7846 => 0, 7847 => 0, 7848 => 0, 7849 => 0, 7850 => 0, 7851 => 0, 7852 => 0, 7853 => 0, 7854 => 0, 7855 => 0, 7856 => 0, 7857 => 1, 7858 => 1, 7859 => 1, 7860 => 1, 7861 => 1, 7862 => 1, 7863 => 1, 7864 => 1, 7865 => 1, 7866 => 1, 7867 => 1, 7868 => 0, 7869 => 0, 7870 => 0, 7871 => 0, 7872 => 0, 7873 => 0, 7874 => 0, 7875 => 0, 7876 => 0, 7877 => 0, 7878 => 0, 7879 => 0, 7880 => 0, 7881 => 0, 7882 => 0, 7883 => 1, 7884 => 1, 7885 => 1, 7886 => 1, 7887 => 1, 7888 => 1, 7889 => 1, 7890 => 1, 7891 => 1, 7892 => 1, 7893 => 1, 7894 => 1, 7895 => 1, 7896 => 1, 7897 => 1, 
7898 => 1, 7899 => 1, 7900 => 1, 7901 => 1, 7902 => 1, 7903 => 1, 7904 => 1, 7905 => 1, 7906 => 1, 7907 => 1, 7908 => 1, 7909 => 1, 7910 => 1, 7911 => 
1, 7912 => 1, 7913 => 0, 7914 => 0, 7915 => 0, 7916 => 0, 7917 => 0, 7918 => 0, 7919 => 0, 7920 => 0, 7921 => 1, 7922 => 1, 7923 => 1, 7924 => 1, 7925 
=> 1, 7926 => 1, 7927 => 1, 7928 => 1, 7929 => 1, 7930 => 1, 7931 => 1, 7932 => 0, 7933 => 0, 7934 => 0, 7935 => 0, 7936 => 0, 7937 => 0, 7938 => 0, 7939 => 0, 7940 => 0, 7941 => 0, 7942 => 0, 7943 => 0, 7944 => 0, 7945 => 0, 7946 => 0, 7947 => 0, 7948 => 0, 7949 => 0, 7950 => 0, 7951 => 0, 7952 => 0, 7953 => 0, 7954 => 0, 7955 => 0, 7956 => 0, 7957 => 0, 7958 => 0, 7959 => 0, 7960 => 0, 7961 => 0, 7962 => 0, 7963 => 0, 7964 => 0, 7965 => 0, 7966 => 0, 7967 => 0, 7968 => 0, 7969 => 0, 7970 => 0, 7971 => 0, 7972 => 0, 7973 => 0, 7974 => 0, 7975 => 0, 7976 => 0, 7977 => 0, 7978 => 1, 7979 => 1, 7980 => 1, 7981 => 1, 7982 => 1, 7983 => 1, 7984 => 1, 7985 => 1, 7986 => 1, 7987 => 1, 7988 => 1, 7989 => 1, 7990 => 1, 7991 => 1, 7992 => 1, 7993 => 1, 7994 => 1, 7995 => 1, 7996 => 1, 7997 => 1, 7998 => 1, 7999 => 1, 8000 => 1, 8001 => 1, 8002 => 1, 8003 => 1, 8004 => 1, 8005 => 1, 8006 => 1, 8007 => 1, 8008 => 1, 8009 => 0, 8010 => 0, 8011 => 0, 8012 => 0, 8013 => 0, 8014 => 0, 8015 => 0, 8016 => 0, 8017 => 0, 8018 => 0, 8019 => 0, 8020 => 0, 8021 => 0, 8022 => 0, 8023 => 1, 8024 => 1, 8025 => 1, 8026 => 1, 8027 => 1, 8028 => 1, 8029 => 1, 8030 => 1, 8031 => 1, 8032 => 1, 8033 => 1, 8034 => 0, 8035 => 0, 8036 => 0, 8037 => 0, 8038 => 0, 8039 => 0, 8040 => 0, 8041 => 0, 8042 => 0, 8043 => 0, 8044 => 0, 8045 => 0, 8046 => 0, 8047 => 0, 8048 => 0, 
8049 => 0, 8050 => 0, 8051 => 0, 8052 => 0, 8053 => 0, 8054 => 0, 8055 => 1, 8056 => 1, 8057 => 1, 8058 => 1, 8059 => 1, 8060 => 1, 8061 => 1, 8062 => 
1, 8063 => 1, 8064 => 1, 8065 => 1, 8066 => 0, 8067 => 0, 8068 => 0, 8069 => 0, 8070 => 0, 8071 => 0, 8072 => 0, 8073 => 0, 8074 => 0, 8075 => 0, 8076 
=> 0, 8077 => 0, 8078 => 0, 8079 => 0, 8080 => 0, 8081 => 1, 8082 => 1, 8083 => 1, 8084 => 1, 8085 => 1, 8086 => 1, 8087 => 1, 8088 => 1, 8089 => 1, 8090 => 1, 8091 => 1, 8092 => 1, 8093 => 1, 8094 => 1, 8095 => 1, 8096 => 1, 8097 => 1, 8098 => 1, 8099 => 1, 8100 => 1, 8101 => 1, 8102 => 1, 8103 => 1, 8104 => 1, 8105 => 1, 8106 => 1, 8107 => 1, 8108 => 1, 8109 => 1, 8110 => 1, 8111 => 0, 8112 => 0, 8113 => 0, 8114 => 0, 8115 => 0, 8116 => 0, 8117 => 0, 8118 => 0, 8119 => 1, 8120 => 1, 8121 => 1, 8122 => 1, 8123 => 1, 8124 => 1, 8125 => 1, 8126 => 1, 8127 => 1, 8128 => 1, 8129 => 1, 8130 => 0, 8131 => 0, 8132 => 0, 8133 => 0, 8134 => 0, 8135 => 0, 8136 => 0, 8137 => 0, 8138 => 0, 8139 => 0, 8140 => 0, 8141 => 0, 8142 => 0, 8143 => 0, 8144 => 0, 8145 => 0, 8146 => 0, 8147 => 0, 8148 => 0, 8149 => 0, 8150 => 0, 8151 => 0, 8152 => 0, 8153 => 0, 8154 => 0, 8155 => 0, 8156 => 0, 8157 => 0, 8158 => 0, 8159 => 0, 8160 => 0, 8161 => 0, 8162 => 0, 8163 => 0, 8164 => 0, 8165 => 0, 8166 => 0, 8167 => 0, 8168 => 0, 8169 => 0, 8170 => 0, 8171 => 0, 8172 => 0, 8173 => 0, 8174 => 0, 8175 => 0, 8176 => 1, 8177 => 1, 8178 => 1, 8179 => 1, 8180 => 1, 8181 => 1, 8182 => 1, 8183 => 1, 8184 => 1, 8185 => 1, 8186 => 1, 8187 => 1, 8188 => 1, 8189 => 1, 8190 => 1, 8191 => 1, 8192 => 1, 8193 => 1, 8194 => 1, 8195 => 1, 8196 => 1, 8197 => 1, 8198 => 1, 8199 => 1, 
8200 => 1, 8201 => 1, 8202 => 1, 8203 => 1, 8204 => 1, 8205 => 1, 8206 => 1, 8207 => 0, 8208 => 0, 8209 => 0, 8210 => 0, 8211 => 0, 8212 => 0, 8213 => 
0, 8214 => 0, 8215 => 0, 8216 => 0, 8217 => 0, 8218 => 0, 8219 => 0, 8220 => 0, 8221 => 1, 8222 => 1, 8223 => 1, 8224 => 1, 8225 => 1, 8226 => 1, 8227 
=> 1, 8228 => 1, 8229 => 1, 8230 => 1, 8231 => 1, 8232 => 0, 8233 => 0, 8234 => 0, 8235 => 0, 8236 => 0, 8237 => 0, 8238 => 0, 8239 => 0, 8240 => 0, 8241 => 0, 8242 => 0, 8243 => 0, 8244 => 0, 8245 => 0, 8246 => 0, 8247 => 0, 8248 => 0, 8249 => 0, 8250 => 0, 8251 => 0, 8252 => 0, 8253 => 1, 8254 => 1, 8255 => 1, 8256 => 1, 8257 => 1, 8258 => 1, 8259 => 1, 8260 => 1, 8261 => 1, 8262 => 1, 8263 => 1, 8264 => 0, 8265 => 0, 8266 => 0, 8267 => 0, 8268 => 0, 8269 => 0, 8270 => 0, 8271 => 0, 8272 => 0, 8273 => 0, 8274 => 0, 8275 => 0, 8276 => 0, 8277 => 0, 8278 => 0, 8279 => 1, 8280 => 1, 8281 => 1, 8282 => 1, 8283 => 1, 8284 => 1, 8285 => 1, 8286 => 1, 8287 => 1, 8288 => 1, 8289 => 1, 8290 => 1, 8291 => 1, 8292 => 1, 8293 => 1, 8294 => 1, 8295 => 1, 8296 => 1, 8297 => 1, 8298 => 1, 8299 => 1, 8300 => 1, 8301 => 1, 8302 => 1, 8303 => 1, 8304 => 1, 8305 => 1, 8306 => 1, 8307 => 1, 8308 => 1, 8309 => 0, 8310 => 0, 8311 => 0, 8312 => 0, 8313 => 0, 8314 => 0, 8315 => 0, 8316 => 0, 8317 => 1, 8318 => 1, 8319 => 1, 8320 => 1, 8321 => 1, 8322 => 1, 8323 => 1, 8324 => 1, 8325 => 1, 8326 => 1, 8327 => 1, 8328 => 0, 8329 => 0, 8330 => 0, 8331 => 0, 8332 => 0, 8333 => 0, 8334 => 0, 8335 => 0, 8336 => 0, 8337 => 0, 8338 => 0, 8339 => 0, 8340 => 0, 8341 => 0, 8342 => 0, 8343 => 0, 8344 => 0, 8345 => 0, 8346 => 0, 8347 => 0, 8348 => 0, 8349 => 0, 8350 => 0, 
8351 => 0, 8352 => 0, 8353 => 0, 8354 => 0, 8355 => 0, 8356 => 0, 8357 => 0, 8358 => 0, 8359 => 0, 8360 => 0, 8361 => 0, 8362 => 0, 8363 => 0, 8364 => 
0, 8365 => 0, 8366 => 0, 8367 => 0, 8368 => 0, 8369 => 0, 8370 => 0, 8371 => 0, 8372 => 0, 8373 => 0, 8374 => 1, 8375 => 1, 8376 => 1, 8377 => 1, 8378 
=> 1, 8379 => 1, 8380 => 1, 8381 => 1, 8382 => 1, 8383 => 1, 8384 => 1, 8385 => 1, 8386 => 1, 8387 => 1, 8388 => 1, 8389 => 1, 8390 => 1, 8391 => 1, 8392 => 1, 8393 => 1, 8394 => 1, 8395 => 1, 8396 => 1, 8397 => 1, 8398 => 1, 8399 => 1, 8400 => 1, 8401 => 1, 8402 => 1, 8403 => 1, 8404 => 1, 8405 => 0, 8406 => 0, 8407 => 0, 8408 => 0, 8409 => 0, 8410 => 0, 8411 => 0, 8412 => 0, 8413 => 0, 8414 => 0, 8415 => 0, 8416 => 0, 8417 => 0, 8418 => 0, 8419 => 1, 8420 => 1, 8421 => 1, 8422 => 1, 8423 => 1, 8424 => 1, 8425 => 1, 8426 => 1, 8427 => 1, 8428 => 1, 8429 => 1, 8430 => 0, 8431 => 0, 8432 => 0, 8433 => 0, 8434 => 0, 8435 => 0, 8436 => 0, 8437 => 0, 8438 => 0, 8439 => 0, 8440 => 0, 8441 => 0, 8442 => 0, 8443 => 0, 8444 => 0, 8445 => 0, 8446 => 0, 8447 => 0, 8448 => 0, 8449 => 0, 8450 => 0, 8451 => 1, 8452 => 1, 8453 => 1, 8454 => 1, 8455 => 1, 8456 => 1, 8457 => 1, 8458 => 1, 8459 => 1, 8460 => 1, 8461 => 1, 8462 => 0, 8463 => 0, 8464 => 0, 8465 => 0, 8466 => 0, 8467 => 0, 8468 => 0, 8469 => 0, 8470 => 0, 8471 => 0, 8472 => 0, 8473 => 0, 8474 => 0, 8475 => 0, 8476 => 0, 8477 => 1, 8478 => 1, 8479 => 1, 8480 => 1, 8481 => 1, 8482 => 1, 8483 => 1, 8484 => 1, 8485 => 1, 8486 => 1, 8487 => 1, 8488 => 1, 8489 => 1, 8490 => 1, 8491 => 1, 8492 => 1, 8493 => 1, 8494 => 1, 8495 => 1, 8496 => 1, 8497 => 1, 8498 => 1, 8499 => 1, 8500 => 1, 8501 => 1, 
8502 => 1, 8503 => 1, 8504 => 1, 8505 => 1, 8506 => 1, 8507 => 0, 8508 => 0, 8509 => 0, 8510 => 0, 8511 => 0, 8512 => 0, 8513 => 0, 8514 => 0, 8515 => 
1, 8516 => 1, 8517 => 1, 8518 => 1, 8519 => 1, 8520 => 1, 8521 => 1, 8522 => 1, 8523 => 1, 8524 => 1, 8525 => 1, 8526 => 0, 8527 => 0, 8528 => 0, 8529 
=> 0, 8530 => 0, 8531 => 0, 8532 => 0, 8533 => 0, 8534 => 0, 8535 => 0, 8536 => 0, 8537 => 0, 8538 => 0, 8539 => 0, 8540 => 0, 8541 => 0, 8542 => 0, 8543 => 0, 8544 => 0, 8545 => 0, 8546 => 0, 8547 => 0, 8548 => 0, 8549 => 0, 8550 => 0, 8551 => 0, 8552 => 0, 8553 => 0, 8554 => 0, 8555 => 0, 8556 => 0, 8557 => 0, 8558 => 0, 8559 => 0, 8560 => 0, 8561 => 0, 8562 => 0, 8563 => 0, 8564 => 0, 8565 => 0, 8566 => 0, 8567 => 0, 8568 => 0, 8569 => 0, 8570 => 0, 8571 => 0, 8572 => 1, 8573 => 1, 8574 => 1, 8575 => 1, 8576 => 1, 8577 => 1, 8578 => 1, 8579 => 1, 8580 => 1, 8581 => 1, 8582 => 1, 8583 => 1, 8584 => 1, 8585 => 1, 8586 => 1, 8587 => 1, 8588 => 1, 8589 => 1, 8590 => 1, 8591 => 1, 8592 => 1, 8593 => 1, 8594 => 1, 8595 => 1, 8596 => 1, 8597 => 1, 8598 => 1, 8599 => 1, 8600 => 1, 8601 => 1, 8602 => 1, 8603 => 0, 8604 => 0, 8605 => 0, 8606 => 0, 8607 => 0, 8608 => 0, 8609 => 0, 8610 => 0, 8611 => 0, 8612 => 0, 8613 => 0, 8614 => 0, 8615 => 0, 8616 => 0, 8617 => 1, 8618 => 1, 8619 => 1, 8620 => 1, 8621 => 1, 8622 => 1, 8623 => 1, 8624 => 1, 8625 => 1, 8626 => 1, 8627 => 1, 8628 => 0, 8629 => 0, 8630 => 0, 8631 => 0, 8632 => 0, 8633 => 0, 8634 => 0, 8635 => 0, 8636 => 0, 8637 => 0, 8638 => 0, 8639 => 0, 8640 => 0, 8641 => 0, 8642 => 0, 8643 => 0, 8644 => 0, 8645 => 0, 8646 => 0, 8647 => 0, 8648 => 0, 8649 => 1, 8650 => 1, 8651 => 1, 8652 => 1, 
8653 => 1, 8654 => 1, 8655 => 1, 8656 => 1, 8657 => 1, 8658 => 1, 8659 => 1, 8660 => 0, 8661 => 0, 8662 => 0, 8663 => 0, 8664 => 0, 8665 => 0, 8666 => 
0, 8667 => 0, 8668 => 0, 8669 => 0, 8670 => 0, 8671 => 0, 8672 => 0, 8673 => 0, 8674 => 0, 8675 => 1, 8676 => 1, 8677 => 1, 8678 => 1, 8679 => 1, 8680 
=> 1, 8681 => 1, 8682 => 1, 8683 => 1, 8684 => 1, 8685 => 1, 8686 => 1, 8687 => 1, 8688 => 1, 8689 => 1, 8690 => 1, 8691 => 1, 8692 => 1, 8693 => 1, 8694 => 1, 8695 => 1, 8696 => 1, 8697 => 1, 8698 => 1, 8699 => 1, 8700 => 1, 8701 => 1, 8702 => 1, 8703 => 1, 8704 => 1, 8705 => 0, 8706 => 0, 8707 => 0, 8708 => 0, 8709 => 0, 8710 => 0, 8711 => 0, 8712 => 0, 8713 => 1, 8714 => 1, 8715 => 1, 8716 => 1, 8717 => 1, 8718 => 1, 8719 => 1, 8720 => 1, 8721 => 1, 8722 => 1, 8723 => 1, 8724 => 0, 8725 => 0, 8726 => 0, 8727 => 0, 8728 => 0, 8729 => 0, 8730 => 0, 8731 => 0, 8732 => 0, 8733 => 0, 8734 => 0, 8735 => 0, 8736 => 0, 8737 => 0, 8738 => 0, 8739 => 0, 8740 => 0, 8741 => 0, 8742 => 0, 8743 => 0, 8744 => 0, 8745 => 0, 8746 => 0, 8747 => 0, 8748 => 0, 8749 => 0, 8750 => 0, 8751 => 0, 8752 => 0, 8753 => 0, 8754 => 0, 8755 => 0, 8756 => 0, 8757 => 0, 8758 => 0, 8759 => 0, 8760 => 0, 8761 => 0, 8762 => 0, 8763 => 0, 8764 => 0, 8765 => 0, 8766 => 0, 8767 => 0, 8768 => 0, 8769 => 0, 8770 => 1, 8771 => 1, 8772 => 1, 8773 => 1, 8774 => 1, 8775 => 1, 8776 => 1, 8777 => 1, 8778 => 1, 8779 => 1, 8780 => 1, 8781 => 1, 8782 => 1, 8783 => 1, 8784 => 1, 8785 => 1, 8786 => 1, 8787 => 1, 8788 => 1, 8789 => 1, 8790 => 1, 8791 => 1, 8792 => 1, 8793 => 1, 8794 => 1, 8795 => 1, 8796 => 1, 8797 => 1, 8798 => 1, 8799 => 1, 8800 => 1, 8801 => 0, 8802 => 0, 8803 => 0, 
8804 => 0, 8805 => 0, 8806 => 0, 8807 => 0, 8808 => 0, 8809 => 0, 8810 => 0, 8811 => 0, 8812 => 0, 8813 => 0, 8814 => 0, 8815 => 1, 8816 => 1, 8817 => 
1, 8818 => 1, 8819 => 1, 8820 => 1, 8821 => 1, 8822 => 1, 8823 => 1, 8824 => 1, 8825 => 1, 8826 => 0, 8827 => 0, 8828 => 0, 8829 => 0, 8830 => 0, 8831 
=> 0, 8832 => 0, 8833 => 0, 8834 => 0, 8835 => 0, 8836 => 0, 8837 => 0, 8838 => 0, 8839 => 0, 8840 => 0, 8841 => 0, 8842 => 0, 8843 => 0, 8844 => 0, 8845 => 0, 8846 => 0, 8847 => 1, 8848 => 1, 8849 => 1, 8850 => 1, 8851 => 1, 8852 => 1, 8853 => 1, 8854 => 1, 8855 => 1, 8856 => 1, 8857 => 1, 8858 => 0, 8859 => 0, 8860 => 0, 8861 => 0, 8862 => 0, 8863 => 0, 8864 => 0, 8865 => 0, 8866 => 0, 8867 => 0, 8868 => 0, 8869 => 0, 8870 => 0, 8871 => 0, 8872 => 0, 8873 => 1, 8874 => 1, 8875 => 1, 8876 => 1, 8877 => 1, 8878 => 1, 8879 => 1, 8880 => 1, 8881 => 1, 8882 => 1, 8883 => 1, 8884 => 1, 8885 => 1, 8886 => 1, 8887 => 1, 8888 => 1, 8889 => 1, 8890 => 1, 8891 => 1, 8892 => 1, 8893 => 1, 8894 => 1, 8895 => 1, 8896 => 1, 8897 => 1, 8898 => 1, 8899 => 1, 8900 => 1, 8901 => 1, 8902 => 1, 8903 => 0, 8904 => 0, 8905 => 0, 8906 => 0, 8907 => 0, 8908 => 0, 8909 => 0
	
	);
	constant rom_game: rom_bitmap_title := (
	0 => 0, 1 => 0, 2 => 0, 3 => 0, 4 => 0, 5 => 0, 6 => 0, 7 => 1, 8 => 1, 9 => 1, 10 => 1, 11 => 1, 12 => 1, 13 => 1, 14 => 1, 15 => 1, 16 => 1, 17 => 1, 18 => 1, 19 => 1, 20 => 1, 21 => 1, 22 => 1, 23 => 1, 24 => 1, 25 => 1, 26 => 1, 27 => 1, 28 => 1, 29 => 1, 30 => 1, 31 => 1, 32 => 1, 33 => 1, 34 => 
1, 35 => 1, 36 => 1, 37 => 1, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 0, 45 => 0, 46 => 0, 47 => 0, 48 => 0, 49 => 0, 50 => 0, 51 => 0, 52 => 0, 53 => 0, 54 => 0, 55 => 0, 56 => 0, 57 => 0, 58 => 0, 59 => 0, 60 => 0, 61 => 0, 62 => 0, 63 => 0, 64 => 0, 65 => 1, 66 => 1, 67 => 1, 68 => 1, 69 => 1, 70 => 1, 71 => 1, 72 => 1, 73 => 1, 74 => 1, 75 => 1, 76 => 1, 77 => 1, 78 => 1, 79 => 1, 80 => 1, 81 => 1, 82 => 1, 83 => 0, 84 => 0, 
85 => 0, 86 => 0, 87 => 0, 88 => 0, 89 => 0, 90 => 0, 91 => 0, 92 => 0, 93 => 0, 94 => 0, 95 => 0, 96 => 0, 97 => 0, 98 => 0, 99 => 0, 100 => 0, 101 => 0, 102 => 0, 103 => 0, 104 => 1, 105 => 1, 106 => 1, 107 => 1, 108 => 1, 109 => 0, 110 => 0, 111 => 0, 112 => 0, 113 => 0, 114 => 0, 115 => 0, 116 => 
0, 117 => 0, 118 => 0, 119 => 0, 120 => 0, 121 => 0, 122 => 0, 123 => 0, 124 => 0, 125 => 0, 126 => 0, 127 => 0, 128 => 0, 129 => 0, 130 => 0, 131 => 0, 132 => 0, 133 => 0, 134 => 0, 135 => 0, 136 => 0, 137 => 0, 138 => 0, 139 => 0, 140 => 0, 141 => 0, 142 => 1, 143 => 1, 144 => 1, 145 => 1, 146 => 1, 147 => 0, 148 => 0, 149 => 0, 150 => 0, 151 => 0, 152 => 0, 153 => 0, 154 => 0, 155 => 1, 156 => 1, 157 => 1, 158 => 1, 159 => 1, 160 => 1, 161 => 1, 
162 => 1, 163 => 1, 164 => 1, 165 => 1, 166 => 1, 167 => 1, 168 => 1, 169 => 1, 170 => 1, 171 => 1, 172 => 1, 173 => 1, 174 => 1, 175 => 1, 176 => 1, 177 => 1, 178 => 1, 179 => 1, 180 => 1, 181 => 1, 182 => 1, 183 => 1, 184 => 1, 185 => 1, 186 => 1, 187 => 1, 188 => 1, 189 => 1, 190 => 1, 191 => 1, 192 => 1, 193 => 1, 194 => 1, 195 => 1, 196 => 1, 197 => 1, 198 => 1, 199 => 0, 200 => 0, 201 => 0, 202 => 0, 203 => 0, 204 => 0, 205 => 0, 206 => 0, 207 => 1, 208 => 1, 209 => 1, 210 => 1, 211 => 1, 212 => 1, 213 => 1, 214 => 1, 215 => 1, 216 => 1, 217 => 1, 218 => 1, 219 => 1, 220 => 1, 221 => 1, 222 
=> 1, 223 => 1, 224 => 1, 225 => 1, 226 => 1, 227 => 1, 228 => 1, 229 => 1, 230 => 1, 231 => 1, 232 => 1, 233 => 1, 234 => 1, 235 => 1, 236 => 1, 237 => 1, 238 => 0, 239 => 0, 240 => 0, 241 => 0, 242 => 0, 243 => 0, 244 => 0, 245 => 0, 246 => 0, 247 => 0, 248 => 0, 249 => 0, 250 => 0, 251 => 0, 252 => 0, 253 => 0, 254 => 0, 255 => 0, 256 => 0, 257 => 0, 258 => 0, 259 => 0, 260 => 0, 261 => 0, 262 => 0, 263 => 0, 264 => 0, 265 => 1, 266 => 1, 267 => 
1, 268 => 1, 269 => 1, 270 => 1, 271 => 1, 272 => 1, 273 => 1, 274 => 1, 275 => 1, 276 => 1, 277 => 1, 278 => 1, 279 => 1, 280 => 1, 281 => 1, 282 => 1, 283 => 0, 284 => 0, 285 => 0, 286 => 0, 287 => 0, 288 => 0, 289 => 0, 290 => 0, 291 => 0, 292 => 0, 293 => 0, 294 => 0, 295 => 0, 296 => 0, 297 => 0, 298 => 0, 299 => 0, 300 => 0, 301 => 0, 302 => 0, 303 => 0, 304 => 1, 305 => 1, 306 => 1, 307 => 1, 308 => 1, 309 => 0, 310 => 0, 311 => 0, 312 => 0, 
313 => 0, 314 => 0, 315 => 0, 316 => 0, 317 => 0, 318 => 0, 319 => 0, 320 => 0, 321 => 0, 322 => 0, 323 => 0, 324 => 0, 325 => 0, 326 => 0, 327 => 0, 328 => 0, 329 => 0, 330 => 0, 331 => 0, 332 => 0, 333 => 0, 334 => 0, 335 => 0, 336 => 0, 337 => 0, 338 => 0, 339 => 0, 340 => 0, 341 => 0, 342 => 1, 343 => 1, 344 => 1, 345 => 1, 346 => 1, 347 => 0, 348 => 0, 349 => 0, 350 => 0, 351 => 0, 352 => 0, 353 => 0, 354 => 0, 355 => 1, 356 => 1, 357 => 1, 358 => 1, 359 => 1, 360 => 1, 361 => 1, 362 => 1, 363 => 1, 364 => 1, 365 => 1, 366 => 1, 367 => 1, 368 => 1, 369 => 1, 370 => 1, 371 => 1, 372 => 1, 373 
=> 1, 374 => 1, 375 => 1, 376 => 1, 377 => 1, 378 => 1, 379 => 1, 380 => 1, 381 => 1, 382 => 1, 383 => 1, 384 => 1, 385 => 1, 386 => 1, 387 => 1, 388 => 1, 389 => 1, 390 => 1, 391 => 1, 392 => 1, 393 => 1, 394 => 1, 395 => 1, 396 => 1, 397 => 1, 398 => 1, 399 => 0, 400 => 0, 401 => 0, 402 => 0, 403 => 0, 404 => 0, 405 => 0, 406 => 0, 407 => 1, 408 => 1, 409 => 1, 410 => 1, 411 => 1, 412 => 1, 413 => 1, 414 => 1, 415 => 1, 416 => 1, 417 => 1, 418 => 
1, 419 => 1, 420 => 1, 421 => 1, 422 => 1, 423 => 1, 424 => 1, 425 => 1, 426 => 1, 427 => 1, 428 => 1, 429 => 1, 430 => 1, 431 => 1, 432 => 1, 433 => 1, 434 => 1, 435 => 1, 436 => 1, 437 => 1, 438 => 0, 439 => 0, 440 => 0, 441 => 0, 442 => 0, 443 => 0, 444 => 0, 445 => 0, 446 => 0, 447 => 0, 448 => 0, 449 => 0, 450 => 0, 451 => 0, 452 => 0, 453 => 0, 454 => 0, 455 => 0, 456 => 0, 457 => 0, 458 => 0, 459 => 0, 460 => 0, 461 => 0, 462 => 0, 463 => 0, 
464 => 0, 465 => 1, 466 => 1, 467 => 1, 468 => 1, 469 => 1, 470 => 1, 471 => 1, 472 => 1, 473 => 1, 474 => 1, 475 => 1, 476 => 1, 477 => 1, 478 => 1, 479 => 1, 480 => 1, 481 => 1, 482 => 1, 483 => 0, 484 => 0, 485 => 0, 486 => 0, 487 => 0, 488 => 0, 489 => 0, 490 => 0, 491 => 0, 492 => 0, 493 => 0, 494 => 0, 495 => 0, 496 => 0, 497 => 0, 498 => 0, 499 => 0, 500 => 0, 501 => 0, 502 => 0, 503 => 0, 504 => 1, 505 => 1, 506 => 1, 507 => 1, 508 => 1, 509 => 0, 510 => 0, 511 => 0, 512 => 0, 513 => 0, 514 => 0, 515 => 0, 516 => 0, 517 => 0, 518 => 0, 519 => 0, 520 => 0, 521 => 0, 522 => 0, 523 => 0, 524 
=> 0, 525 => 0, 526 => 0, 527 => 0, 528 => 0, 529 => 0, 530 => 0, 531 => 0, 532 => 0, 533 => 0, 534 => 0, 535 => 0, 536 => 0, 537 => 0, 538 => 0, 539 => 0, 540 => 0, 541 => 0, 542 => 1, 543 => 1, 544 => 1, 545 => 1, 546 => 1, 547 => 0, 548 => 0, 549 => 0, 550 => 0, 551 => 0, 552 => 0, 553 => 0, 554 => 0, 555 => 1, 556 => 1, 557 => 1, 558 => 1, 559 => 1, 560 => 1, 561 => 1, 562 => 1, 563 => 1, 564 => 1, 565 => 1, 566 => 1, 567 => 1, 568 => 1, 569 => 
1, 570 => 1, 571 => 1, 572 => 1, 573 => 1, 574 => 1, 575 => 1, 576 => 1, 577 => 1, 578 => 1, 579 => 1, 580 => 1, 581 => 1, 582 => 1, 583 => 1, 584 => 1, 585 => 1, 586 => 1, 587 => 1, 588 => 1, 589 => 1, 590 => 1, 591 => 1, 592 => 1, 593 => 1, 594 => 1, 595 => 1, 596 => 1, 597 => 1, 598 => 1, 599 => 0, 600 => 0, 601 => 0, 602 => 0, 603 => 0, 604 => 0, 605 => 0, 606 => 0, 607 => 1, 608 => 1, 609 => 1, 610 => 1, 611 => 1, 612 => 1, 613 => 1, 614 => 1, 
615 => 1, 616 => 1, 617 => 1, 618 => 1, 619 => 1, 620 => 1, 621 => 1, 622 => 1, 623 => 1, 624 => 1, 625 => 1, 626 => 1, 627 => 1, 628 => 1, 629 => 1, 630 => 1, 631 => 1, 632 => 1, 633 => 1, 634 => 1, 635 => 1, 636 => 1, 637 => 1, 638 => 0, 639 => 0, 640 => 0, 641 => 0, 642 => 0, 643 => 0, 644 => 0, 645 => 0, 646 => 0, 647 => 0, 648 => 0, 649 => 0, 650 => 0, 651 => 0, 652 => 0, 653 => 0, 654 => 0, 655 => 0, 656 => 0, 657 => 0, 658 => 0, 659 => 0, 660 => 0, 661 => 0, 662 => 0, 663 => 0, 664 => 0, 665 => 1, 666 => 1, 667 => 1, 668 => 1, 669 => 1, 670 => 1, 671 => 1, 672 => 1, 673 => 1, 674 => 1, 675 
=> 1, 676 => 1, 677 => 1, 678 => 1, 679 => 1, 680 => 1, 681 => 1, 682 => 1, 683 => 0, 684 => 0, 685 => 0, 686 => 0, 687 => 0, 688 => 0, 689 => 0, 690 => 0, 691 => 0, 692 => 0, 693 => 0, 694 => 0, 695 => 0, 696 => 0, 697 => 0, 698 => 0, 699 => 0, 700 => 0, 701 => 0, 702 => 0, 703 => 0, 704 => 1, 705 => 1, 706 => 1, 707 => 1, 708 => 1, 709 => 0, 710 => 0, 711 => 0, 712 => 0, 713 => 0, 714 => 0, 715 => 0, 716 => 0, 717 => 0, 718 => 0, 719 => 0, 720 => 
0, 721 => 0, 722 => 0, 723 => 0, 724 => 0, 725 => 0, 726 => 0, 727 => 0, 728 => 0, 729 => 0, 730 => 0, 731 => 0, 732 => 0, 733 => 0, 734 => 0, 735 => 0, 736 => 0, 737 => 0, 738 => 0, 739 => 0, 740 => 0, 741 => 0, 742 => 1, 743 => 1, 744 => 1, 745 => 1, 746 => 1, 747 => 0, 748 => 0, 749 => 0, 750 => 0, 751 => 0, 752 => 0, 753 => 0, 754 => 0, 755 => 1, 756 => 1, 757 => 1, 758 => 1, 759 => 1, 760 => 1, 761 => 1, 762 => 1, 763 => 1, 764 => 1, 765 => 1, 
766 => 1, 767 => 1, 768 => 1, 769 => 1, 770 => 1, 771 => 1, 772 => 1, 773 => 1, 774 => 1, 775 => 1, 776 => 1, 777 => 1, 778 => 1, 779 => 1, 780 => 1, 781 => 1, 782 => 1, 783 => 1, 784 => 1, 785 => 1, 786 => 1, 787 => 1, 788 => 1, 789 => 1, 790 => 1, 791 => 1, 792 => 1, 793 => 1, 794 => 1, 795 => 1, 796 => 1, 797 => 1, 798 => 1, 799 => 0, 800 => 0, 801 => 0, 802 => 0, 803 => 0, 804 => 0, 805 => 0, 806 => 0, 807 => 1, 808 => 1, 809 => 1, 810 => 1, 811 => 1, 812 => 1, 813 => 1, 814 => 1, 815 => 1, 816 => 1, 817 => 1, 818 => 1, 819 => 1, 820 => 1, 821 => 1, 822 => 1, 823 => 1, 824 => 1, 825 => 1, 826 
=> 1, 827 => 1, 828 => 1, 829 => 1, 830 => 1, 831 => 1, 832 => 1, 833 => 1, 834 => 1, 835 => 1, 836 => 1, 837 => 1, 838 => 0, 839 => 0, 840 => 0, 841 => 0, 842 => 0, 843 => 0, 844 => 0, 845 => 0, 846 => 0, 847 => 0, 848 => 0, 849 => 0, 850 => 0, 851 => 0, 852 => 0, 853 => 0, 854 => 0, 855 => 0, 856 => 0, 857 => 0, 858 => 0, 859 => 0, 860 => 0, 861 => 0, 862 => 0, 863 => 0, 864 => 0, 865 => 1, 866 => 1, 867 => 1, 868 => 1, 869 => 1, 870 => 1, 871 => 
1, 872 => 1, 873 => 1, 874 => 1, 875 => 1, 876 => 1, 877 => 1, 878 => 1, 879 => 1, 880 => 1, 881 => 1, 882 => 1, 883 => 0, 884 => 0, 885 => 0, 886 => 0, 887 => 0, 888 => 0, 889 => 0, 890 => 0, 891 => 0, 892 => 0, 893 => 0, 894 => 0, 895 => 0, 896 => 0, 897 => 0, 898 => 0, 899 => 0, 900 => 0, 901 => 0, 902 => 0, 903 => 0, 904 => 1, 905 => 1, 906 => 1, 907 => 1, 908 => 1, 909 => 0, 910 => 0, 911 => 0, 912 => 0, 913 => 0, 914 => 0, 915 => 0, 916 => 0, 
917 => 0, 918 => 0, 919 => 0, 920 => 0, 921 => 0, 922 => 0, 923 => 0, 924 => 0, 925 => 0, 926 => 0, 927 => 0, 928 => 0, 929 => 0, 930 => 0, 931 => 0, 932 => 0, 933 => 0, 934 => 0, 935 => 0, 936 => 0, 937 => 0, 938 => 0, 939 => 0, 940 => 0, 941 => 0, 942 => 1, 943 => 1, 944 => 1, 945 => 1, 946 => 1, 947 => 0, 948 => 0, 949 => 0, 950 => 0, 951 => 0, 952 => 0, 953 => 0, 954 => 0, 955 => 1, 956 => 1, 957 => 1, 958 => 1, 959 => 1, 960 => 1, 961 => 1, 962 => 1, 963 => 1, 964 => 1, 965 => 1, 966 => 1, 967 => 1, 968 => 1, 969 => 1, 970 => 1, 971 => 1, 972 => 1, 973 => 1, 974 => 1, 975 => 1, 976 => 1, 977 
=> 1, 978 => 1, 979 => 1, 980 => 1, 981 => 1, 982 => 1, 983 => 1, 984 => 1, 985 => 1, 986 => 1, 987 => 1, 988 => 1, 989 => 1, 990 => 1, 991 => 1, 992 => 1, 993 => 1, 994 => 1, 995 => 1, 996 => 1, 997 => 1, 998 => 1, 999 => 0, 1000 => 0, 1001 => 0, 1002 => 0, 1003 => 0, 1004 => 0, 1005 => 0, 1006 => 0, 1007 => 1, 1008 => 1, 1009 => 1, 1010 => 1, 1011 => 1, 1012 => 1, 1013 => 1, 1014 => 1, 1015 => 1, 1016 => 1, 1017 => 1, 1018 => 1, 1019 => 1, 1020 => 1, 1021 => 1, 1022 => 1, 1023 => 1, 1024 => 1, 1025 => 1, 1026 => 1, 1027 => 1, 1028 => 1, 1029 => 1, 1030 => 1, 1031 => 1, 1032 => 1, 1033 => 1, 1034 => 1, 1035 => 1, 1036 => 1, 1037 => 1, 1038 => 0, 1039 => 0, 1040 => 0, 1041 => 0, 1042 => 0, 1043 => 0, 1044 => 0, 1045 => 0, 1046 => 0, 1047 => 0, 1048 => 0, 1049 => 0, 1050 => 0, 1051 => 0, 1052 => 0, 1053 => 0, 1054 => 0, 1055 => 0, 1056 => 0, 1057 => 0, 1058 => 0, 1059 => 0, 1060 => 0, 1061 => 0, 1062 => 0, 1063 => 0, 1064 => 0, 1065 => 1, 1066 => 1, 1067 => 1, 1068 => 1, 1069 => 1, 1070 => 1, 1071 => 1, 1072 => 1, 1073 => 1, 1074 => 1, 1075 => 1, 1076 => 1, 1077 => 1, 1078 => 1, 1079 => 1, 1080 => 1, 1081 => 1, 1082 => 1, 1083 => 0, 1084 => 0, 1085 => 0, 1086 => 0, 1087 => 0, 1088 => 0, 1089 => 0, 1090 => 0, 1091 => 0, 1092 => 0, 1093 => 0, 1094 => 0, 1095 => 0, 1096 => 0, 1097 => 0, 1098 => 0, 1099 => 0, 1100 => 0, 1101 => 0, 1102 => 0, 
1103 => 0, 1104 => 1, 1105 => 1, 1106 => 1, 1107 => 1, 1108 => 1, 1109 => 0, 1110 => 0, 1111 => 0, 1112 => 0, 1113 => 0, 1114 => 0, 1115 => 0, 1116 => 
0, 1117 => 0, 1118 => 0, 1119 => 0, 1120 => 0, 1121 => 0, 1122 => 0, 1123 => 0, 1124 => 0, 1125 => 0, 1126 => 0, 1127 => 0, 1128 => 0, 1129 => 0, 1130 
=> 0, 1131 => 0, 1132 => 0, 1133 => 0, 1134 => 0, 1135 => 0, 1136 => 0, 1137 => 0, 1138 => 0, 1139 => 0, 1140 => 0, 1141 => 0, 1142 => 1, 1143 => 1, 1144 => 1, 1145 => 1, 1146 => 1, 1147 => 0, 1148 => 0, 1149 => 0, 1150 => 0, 1151 => 0, 1152 => 0, 1153 => 0, 1154 => 0, 1155 => 1, 1156 => 1, 1157 => 1, 1158 => 1, 1159 => 1, 1160 => 1, 1161 => 1, 1162 => 1, 1163 => 1, 1164 => 1, 1165 => 1, 1166 => 1, 1167 => 1, 1168 => 1, 1169 => 1, 1170 => 1, 1171 => 1, 1172 => 1, 1173 => 1, 1174 => 1, 1175 => 1, 1176 => 1, 1177 => 1, 1178 => 1, 1179 => 1, 1180 => 1, 1181 => 1, 1182 => 1, 1183 => 1, 1184 => 1, 1185 => 1, 1186 => 1, 1187 => 1, 1188 => 1, 1189 => 1, 1190 => 1, 1191 => 1, 1192 => 1, 1193 => 1, 1194 => 1, 1195 => 1, 1196 => 1, 1197 => 1, 1198 => 1, 1199 => 0, 1200 => 0, 1201 => 0, 1202 => 0, 1203 => 0, 1204 => 0, 1205 => 0, 1206 => 0, 1207 => 1, 1208 => 1, 1209 => 1, 1210 => 1, 1211 => 1, 1212 => 0, 1213 => 0, 1214 => 0, 1215 => 0, 1216 => 0, 1217 => 0, 1218 => 0, 1219 => 0, 1220 => 0, 1221 => 0, 1222 => 0, 1223 => 0, 1224 => 0, 1225 => 0, 1226 => 0, 1227 => 0, 1228 => 0, 1229 => 0, 1230 => 0, 1231 => 0, 1232 => 0, 1233 => 1, 1234 => 1, 1235 => 1, 1236 => 1, 1237 => 1, 1238 => 0, 1239 => 0, 1240 => 0, 1241 => 0, 1242 => 0, 1243 => 0, 1244 => 0, 1245 => 0, 1246 => 0, 1247 => 0, 1248 => 0, 1249 => 0, 1250 => 0, 1251 => 0, 1252 => 0, 1253 => 0, 
1254 => 0, 1255 => 0, 1256 => 0, 1257 => 0, 1258 => 0, 1259 => 0, 1260 => 0, 1261 => 0, 1262 => 0, 1263 => 0, 1264 => 0, 1265 => 1, 1266 => 1, 1267 => 
1, 1268 => 1, 1269 => 1, 1270 => 0, 1271 => 0, 1272 => 0, 1273 => 0, 1274 => 0, 1275 => 0, 1276 => 0, 1277 => 0, 1278 => 1, 1279 => 1, 1280 => 1, 1281 
=> 1, 1282 => 1, 1283 => 0, 1284 => 0, 1285 => 0, 1286 => 0, 1287 => 0, 1288 => 0, 1289 => 0, 1290 => 0, 1291 => 0, 1292 => 0, 1293 => 0, 1294 => 0, 1295 => 0, 1296 => 0, 1297 => 0, 1298 => 0, 1299 => 0, 1300 => 0, 1301 => 0, 1302 => 0, 1303 => 0, 1304 => 1, 1305 => 1, 1306 => 1, 1307 => 1, 1308 => 1, 1309 => 0, 1310 => 0, 1311 => 0, 1312 => 0, 1313 => 0, 1314 => 0, 1315 => 0, 1316 => 0, 1317 => 0, 1318 => 0, 1319 => 0, 1320 => 0, 1321 => 0, 1322 => 0, 1323 => 0, 1324 => 0, 1325 => 0, 1326 => 0, 1327 => 0, 1328 => 0, 1329 => 0, 1330 => 0, 1331 => 0, 1332 => 0, 1333 => 0, 1334 => 0, 1335 => 0, 1336 => 0, 1337 => 0, 1338 => 0, 1339 => 0, 1340 => 0, 1341 => 0, 1342 => 1, 1343 => 1, 1344 => 1, 1345 => 1, 1346 => 1, 1347 => 0, 1348 => 0, 1349 => 0, 1350 => 0, 1351 => 0, 1352 => 0, 1353 => 0, 1354 => 0, 1355 => 1, 1356 => 1, 1357 => 1, 1358 => 1, 1359 => 1, 1360 => 1, 1361 => 1, 1362 => 1, 1363 => 1, 1364 => 1, 1365 => 1, 1366 => 1, 1367 => 0, 1368 => 0, 1369 => 0, 1370 => 0, 1371 => 0, 1372 => 0, 1373 => 0, 1374 => 0, 1375 => 0, 1376 => 0, 1377 => 0, 1378 => 0, 1379 => 0, 1380 => 0, 1381 => 0, 1382 => 0, 1383 => 0, 1384 => 0, 1385 => 0, 1386 => 0, 1387 => 0, 1388 => 0, 1389 => 0, 1390 => 0, 1391 => 0, 1392 => 0, 1393 => 0, 1394 => 0, 1395 => 0, 1396 => 0, 1397 => 0, 1398 => 0, 1399 => 0, 1400 => 0, 1401 => 1, 1402 => 1, 1403 => 1, 1404 => 1, 
1405 => 1, 1406 => 1, 1407 => 1, 1408 => 1, 1409 => 1, 1410 => 1, 1411 => 1, 1412 => 0, 1413 => 0, 1414 => 0, 1415 => 0, 1416 => 0, 1417 => 0, 1418 => 
0, 1419 => 0, 1420 => 0, 1421 => 0, 1422 => 0, 1423 => 0, 1424 => 0, 1425 => 0, 1426 => 0, 1427 => 0, 1428 => 0, 1429 => 0, 1430 => 0, 1431 => 0, 1432 
=> 0, 1433 => 1, 1434 => 1, 1435 => 1, 1436 => 1, 1437 => 1, 1438 => 1, 1439 => 1, 1440 => 1, 1441 => 1, 1442 => 1, 1443 => 1, 1444 => 0, 1445 => 0, 1446 => 0, 1447 => 0, 1448 => 0, 1449 => 0, 1450 => 0, 1451 => 0, 1452 => 0, 1453 => 0, 1454 => 0, 1455 => 0, 1456 => 0, 1457 => 0, 1458 => 0, 1459 => 1, 1460 => 1, 1461 => 1, 1462 => 1, 1463 => 1, 1464 => 1, 1465 => 1, 1466 => 1, 1467 => 1, 1468 => 1, 1469 => 1, 1470 => 0, 1471 => 0, 1472 => 0, 1473 => 0, 1474 => 0, 1475 => 0, 1476 => 0, 1477 => 0, 1478 => 1, 1479 => 1, 1480 => 1, 1481 => 1, 1482 => 1, 1483 => 1, 1484 => 1, 1485 => 1, 1486 => 1, 1487 => 1, 1488 => 1, 1489 => 0, 1490 => 0, 1491 => 0, 1492 => 0, 1493 => 0, 1494 => 0, 1495 => 0, 1496 => 0, 1497 => 0, 1498 => 0, 1499 => 0, 1500 => 0, 1501 => 0, 1502 => 0, 1503 => 0, 1504 => 1, 1505 => 1, 1506 => 1, 1507 => 1, 1508 => 1, 1509 => 1, 1510 => 1, 1511 => 1, 1512 => 1, 1513 => 1, 1514 => 1, 1515 => 1, 1516 => 0, 1517 => 0, 1518 => 0, 1519 => 0, 1520 => 0, 1521 => 0, 1522 => 0, 1523 => 0, 1524 => 0, 1525 => 0, 1526 => 0, 1527 => 0, 1528 => 0, 1529 => 0, 1530 => 0, 1531 => 0, 1532 => 0, 1533 => 0, 1534 => 0, 1535 => 0, 1536 => 1, 1537 => 1, 1538 => 1, 1539 => 1, 1540 => 1, 1541 => 1, 1542 => 1, 1543 => 1, 1544 => 1, 1545 => 1, 1546 => 1, 1547 => 0, 1548 => 0, 1549 => 0, 1550 => 0, 1551 => 0, 1552 => 0, 1553 => 0, 1554 => 0, 1555 => 1, 
1556 => 1, 1557 => 1, 1558 => 1, 1559 => 1, 1560 => 1, 1561 => 1, 1562 => 1, 1563 => 1, 1564 => 1, 1565 => 1, 1566 => 1, 1567 => 0, 1568 => 0, 1569 => 
0, 1570 => 0, 1571 => 0, 1572 => 0, 1573 => 0, 1574 => 0, 1575 => 0, 1576 => 0, 1577 => 0, 1578 => 0, 1579 => 0, 1580 => 0, 1581 => 0, 1582 => 0, 1583 
=> 0, 1584 => 0, 1585 => 0, 1586 => 0, 1587 => 0, 1588 => 0, 1589 => 0, 1590 => 0, 1591 => 0, 1592 => 0, 1593 => 0, 1594 => 0, 1595 => 0, 1596 => 0, 1597 => 0, 1598 => 0, 1599 => 0, 1600 => 0, 1601 => 1, 1602 => 1, 1603 => 1, 1604 => 1, 1605 => 1, 1606 => 1, 1607 => 1, 1608 => 1, 1609 => 1, 1610 => 1, 1611 => 1, 1612 => 0, 1613 => 0, 1614 => 0, 1615 => 0, 1616 => 0, 1617 => 0, 1618 => 0, 1619 => 0, 1620 => 0, 1621 => 0, 1622 => 0, 1623 => 0, 1624 => 0, 1625 => 0, 1626 => 0, 1627 => 0, 1628 => 0, 1629 => 0, 1630 => 0, 1631 => 0, 1632 => 0, 1633 => 1, 1634 => 1, 1635 => 1, 1636 => 1, 1637 => 1, 1638 => 1, 1639 => 1, 1640 => 1, 1641 => 1, 1642 => 1, 1643 => 1, 1644 => 0, 1645 => 0, 1646 => 0, 1647 => 0, 1648 => 0, 1649 => 0, 1650 => 0, 1651 => 0, 1652 => 0, 1653 => 0, 1654 => 0, 1655 => 0, 1656 => 0, 1657 => 0, 1658 => 0, 1659 => 1, 1660 => 1, 1661 => 1, 1662 => 1, 1663 => 1, 1664 => 1, 1665 => 1, 1666 => 1, 1667 => 1, 1668 => 1, 1669 => 1, 1670 => 0, 1671 => 0, 1672 => 0, 1673 => 0, 1674 => 0, 1675 => 0, 1676 => 0, 1677 => 0, 1678 => 1, 1679 => 1, 1680 => 1, 1681 => 1, 1682 => 1, 1683 => 1, 1684 => 1, 1685 => 1, 1686 => 1, 1687 => 1, 1688 => 1, 1689 => 0, 1690 => 0, 1691 => 0, 1692 => 0, 1693 => 0, 1694 => 0, 1695 => 0, 1696 => 0, 1697 => 0, 1698 => 0, 1699 => 0, 1700 => 0, 1701 => 0, 1702 => 0, 1703 => 0, 1704 => 1, 1705 => 1, 1706 => 1, 
1707 => 1, 1708 => 1, 1709 => 1, 1710 => 1, 1711 => 1, 1712 => 1, 1713 => 1, 1714 => 1, 1715 => 1, 1716 => 0, 1717 => 0, 1718 => 0, 1719 => 0, 1720 => 
0, 1721 => 0, 1722 => 0, 1723 => 0, 1724 => 0, 1725 => 0, 1726 => 0, 1727 => 0, 1728 => 0, 1729 => 0, 1730 => 0, 1731 => 0, 1732 => 0, 1733 => 0, 1734 
=> 0, 1735 => 0, 1736 => 1, 1737 => 1, 1738 => 1, 1739 => 1, 1740 => 1, 1741 => 1, 1742 => 1, 1743 => 1, 1744 => 1, 1745 => 1, 1746 => 1, 1747 => 0, 1748 => 0, 1749 => 0, 1750 => 0, 1751 => 0, 1752 => 0, 1753 => 0, 1754 => 0, 1755 => 1, 1756 => 1, 1757 => 1, 1758 => 1, 1759 => 1, 1760 => 1, 1761 => 1, 1762 => 1, 1763 => 1, 1764 => 1, 1765 => 1, 1766 => 1, 1767 => 0, 1768 => 0, 1769 => 0, 1770 => 0, 1771 => 0, 1772 => 0, 1773 => 0, 1774 => 0, 1775 => 0, 1776 => 0, 1777 => 0, 1778 => 0, 1779 => 0, 1780 => 0, 1781 => 0, 1782 => 0, 1783 => 0, 1784 => 0, 1785 => 0, 1786 => 0, 1787 => 0, 1788 => 0, 1789 => 0, 1790 => 0, 1791 => 0, 1792 => 0, 1793 => 0, 1794 => 0, 1795 => 0, 1796 => 0, 1797 => 0, 1798 => 0, 1799 => 0, 1800 => 0, 1801 => 1, 1802 => 1, 1803 => 1, 1804 => 1, 1805 => 1, 1806 => 1, 1807 => 1, 1808 => 1, 1809 => 1, 1810 => 1, 1811 => 1, 1812 => 0, 1813 => 0, 1814 => 0, 1815 => 0, 1816 => 0, 1817 => 0, 1818 => 0, 1819 => 0, 1820 => 0, 1821 => 0, 1822 => 0, 1823 => 0, 1824 => 0, 1825 => 0, 1826 => 0, 1827 => 0, 1828 => 0, 1829 => 0, 1830 => 0, 1831 => 0, 1832 => 0, 1833 => 1, 1834 => 1, 1835 => 1, 1836 => 1, 1837 => 1, 1838 => 1, 1839 => 1, 1840 => 1, 1841 => 1, 1842 => 1, 1843 => 1, 1844 => 0, 1845 => 0, 1846 => 0, 1847 => 0, 1848 => 0, 1849 => 0, 1850 => 0, 1851 => 0, 1852 => 0, 1853 => 0, 1854 => 0, 1855 => 0, 1856 => 0, 1857 => 0, 
1858 => 0, 1859 => 1, 1860 => 1, 1861 => 1, 1862 => 1, 1863 => 1, 1864 => 1, 1865 => 1, 1866 => 1, 1867 => 1, 1868 => 1, 1869 => 1, 1870 => 0, 1871 => 
0, 1872 => 0, 1873 => 0, 1874 => 0, 1875 => 0, 1876 => 0, 1877 => 0, 1878 => 1, 1879 => 1, 1880 => 1, 1881 => 1, 1882 => 1, 1883 => 1, 1884 => 1, 1885 
=> 1, 1886 => 1, 1887 => 1, 1888 => 1, 1889 => 0, 1890 => 0, 1891 => 0, 1892 => 0, 1893 => 0, 1894 => 0, 1895 => 0, 1896 => 0, 1897 => 0, 1898 => 0, 1899 => 0, 1900 => 0, 1901 => 0, 1902 => 0, 1903 => 0, 1904 => 1, 1905 => 1, 1906 => 1, 1907 => 1, 1908 => 1, 1909 => 1, 1910 => 1, 1911 => 1, 1912 => 1, 1913 => 1, 1914 => 1, 1915 => 1, 1916 => 0, 1917 => 0, 1918 => 0, 1919 => 0, 1920 => 0, 1921 => 0, 1922 => 0, 1923 => 0, 1924 => 0, 1925 => 0, 1926 => 0, 1927 => 0, 1928 => 0, 1929 => 0, 1930 => 0, 1931 => 0, 1932 => 0, 1933 => 0, 1934 => 0, 1935 => 0, 1936 => 1, 1937 => 1, 1938 => 1, 1939 => 1, 1940 => 1, 1941 => 1, 1942 => 1, 1943 => 1, 1944 => 1, 1945 => 1, 1946 => 1, 1947 => 0, 1948 => 0, 1949 => 0, 1950 => 0, 1951 => 0, 1952 => 0, 1953 => 0, 1954 => 0, 1955 => 1, 1956 => 1, 1957 => 1, 1958 => 1, 1959 => 1, 1960 => 1, 1961 => 1, 1962 => 1, 1963 => 1, 1964 => 1, 1965 => 1, 1966 => 1, 1967 => 0, 1968 => 0, 1969 => 0, 1970 => 0, 1971 => 0, 1972 => 0, 1973 => 0, 1974 => 0, 1975 => 0, 1976 => 0, 1977 => 0, 1978 => 0, 1979 => 0, 1980 => 0, 1981 => 0, 1982 => 0, 1983 => 0, 1984 => 0, 1985 => 0, 1986 => 0, 1987 => 0, 1988 => 0, 1989 => 0, 1990 => 0, 1991 => 0, 1992 => 0, 1993 => 0, 1994 => 0, 1995 => 0, 1996 => 0, 1997 => 0, 1998 => 0, 1999 => 0, 2000 => 0, 2001 => 1, 2002 => 1, 2003 => 1, 2004 => 1, 2005 => 1, 2006 => 1, 2007 => 1, 2008 => 1, 
2009 => 1, 2010 => 1, 2011 => 1, 2012 => 0, 2013 => 0, 2014 => 0, 2015 => 0, 2016 => 0, 2017 => 0, 2018 => 0, 2019 => 0, 2020 => 0, 2021 => 0, 2022 => 
0, 2023 => 0, 2024 => 0, 2025 => 0, 2026 => 0, 2027 => 0, 2028 => 0, 2029 => 0, 2030 => 0, 2031 => 0, 2032 => 0, 2033 => 1, 2034 => 1, 2035 => 1, 2036 
=> 1, 2037 => 1, 2038 => 1, 2039 => 1, 2040 => 1, 2041 => 1, 2042 => 1, 2043 => 1, 2044 => 0, 2045 => 0, 2046 => 0, 2047 => 0, 2048 => 0, 2049 => 0, 2050 => 0, 2051 => 0, 2052 => 0, 2053 => 0, 2054 => 0, 2055 => 0, 2056 => 0, 2057 => 0, 2058 => 0, 2059 => 1, 2060 => 1, 2061 => 1, 2062 => 1, 2063 => 1, 2064 => 1, 2065 => 1, 2066 => 1, 2067 => 1, 2068 => 1, 2069 => 1, 2070 => 0, 2071 => 0, 2072 => 0, 2073 => 0, 2074 => 0, 2075 => 0, 2076 => 0, 2077 => 0, 2078 => 1, 2079 => 1, 2080 => 1, 2081 => 1, 2082 => 1, 2083 => 1, 2084 => 1, 2085 => 1, 2086 => 1, 2087 => 1, 2088 => 1, 2089 => 0, 2090 => 0, 2091 => 0, 2092 => 0, 2093 => 0, 2094 => 0, 2095 => 0, 2096 => 0, 2097 => 0, 2098 => 0, 2099 => 0, 2100 => 0, 2101 => 0, 2102 => 0, 2103 => 0, 2104 => 1, 2105 => 1, 2106 => 1, 2107 => 1, 2108 => 1, 2109 => 1, 2110 => 1, 2111 => 1, 2112 => 1, 2113 => 1, 2114 => 1, 2115 => 1, 2116 => 0, 2117 => 0, 2118 => 0, 2119 => 0, 2120 => 0, 2121 => 0, 2122 => 0, 2123 => 0, 2124 => 0, 2125 => 0, 2126 => 0, 2127 => 0, 2128 => 0, 2129 => 0, 2130 => 0, 2131 => 0, 2132 => 0, 2133 => 0, 2134 => 0, 2135 => 0, 2136 => 1, 2137 => 1, 2138 => 1, 2139 => 1, 2140 => 1, 2141 => 1, 2142 => 1, 2143 => 1, 2144 => 1, 2145 => 1, 2146 => 1, 2147 => 0, 2148 => 0, 2149 => 0, 2150 => 0, 2151 => 0, 2152 => 0, 2153 => 0, 2154 => 0, 2155 => 1, 2156 => 1, 2157 => 1, 2158 => 1, 2159 => 1, 
2160 => 1, 2161 => 1, 2162 => 1, 2163 => 1, 2164 => 1, 2165 => 1, 2166 => 1, 2167 => 0, 2168 => 0, 2169 => 0, 2170 => 0, 2171 => 0, 2172 => 0, 2173 => 
0, 2174 => 0, 2175 => 0, 2176 => 0, 2177 => 0, 2178 => 0, 2179 => 0, 2180 => 0, 2181 => 0, 2182 => 0, 2183 => 0, 2184 => 0, 2185 => 0, 2186 => 0, 2187 
=> 0, 2188 => 0, 2189 => 0, 2190 => 0, 2191 => 0, 2192 => 0, 2193 => 0, 2194 => 0, 2195 => 0, 2196 => 0, 2197 => 0, 2198 => 0, 2199 => 0, 2200 => 0, 2201 => 1, 2202 => 1, 2203 => 1, 2204 => 1, 2205 => 1, 2206 => 1, 2207 => 1, 2208 => 1, 2209 => 1, 2210 => 1, 2211 => 1, 2212 => 0, 2213 => 0, 2214 => 0, 2215 => 0, 2216 => 0, 2217 => 0, 2218 => 0, 2219 => 0, 2220 => 0, 2221 => 0, 2222 => 0, 2223 => 0, 2224 => 0, 2225 => 0, 2226 => 0, 2227 => 0, 2228 => 0, 2229 => 0, 2230 => 0, 2231 => 0, 2232 => 0, 2233 => 1, 2234 => 1, 2235 => 1, 2236 => 1, 2237 => 1, 2238 => 1, 2239 => 1, 2240 => 1, 2241 => 1, 2242 => 1, 2243 => 1, 2244 => 0, 2245 => 0, 2246 => 0, 2247 => 0, 2248 => 0, 2249 => 0, 2250 => 0, 2251 => 0, 2252 => 0, 2253 => 0, 2254 => 0, 2255 => 0, 2256 => 0, 2257 => 0, 2258 => 0, 2259 => 1, 2260 => 1, 2261 => 1, 2262 => 1, 2263 => 1, 2264 => 1, 2265 => 1, 2266 => 1, 2267 => 1, 2268 => 1, 2269 => 1, 2270 => 0, 2271 => 0, 2272 => 0, 2273 => 0, 2274 => 0, 2275 => 0, 2276 => 0, 2277 => 0, 2278 => 1, 2279 => 1, 2280 => 1, 2281 => 1, 2282 => 1, 2283 => 1, 2284 => 1, 2285 => 1, 2286 => 1, 2287 => 1, 2288 => 1, 2289 => 0, 2290 => 0, 2291 => 0, 2292 => 0, 2293 => 0, 2294 => 0, 2295 => 0, 2296 => 0, 2297 => 0, 2298 => 0, 2299 => 0, 2300 => 0, 2301 => 0, 2302 => 0, 2303 => 0, 2304 => 1, 2305 => 1, 2306 => 1, 2307 => 1, 2308 => 1, 2309 => 1, 2310 => 1, 
2311 => 1, 2312 => 1, 2313 => 1, 2314 => 1, 2315 => 1, 2316 => 0, 2317 => 0, 2318 => 0, 2319 => 0, 2320 => 0, 2321 => 0, 2322 => 0, 2323 => 0, 2324 => 
0, 2325 => 0, 2326 => 0, 2327 => 0, 2328 => 0, 2329 => 0, 2330 => 0, 2331 => 0, 2332 => 0, 2333 => 0, 2334 => 0, 2335 => 0, 2336 => 1, 2337 => 1, 2338 
=> 1, 2339 => 1, 2340 => 1, 2341 => 1, 2342 => 1, 2343 => 1, 2344 => 1, 2345 => 1, 2346 => 1, 2347 => 0, 2348 => 0, 2349 => 0, 2350 => 0, 2351 => 0, 2352 => 0, 2353 => 0, 2354 => 0, 2355 => 1, 2356 => 1, 2357 => 1, 2358 => 1, 2359 => 1, 2360 => 1, 2361 => 1, 2362 => 1, 2363 => 1, 2364 => 1, 2365 => 1, 2366 => 1, 2367 => 0, 2368 => 0, 2369 => 0, 2370 => 0, 2371 => 0, 2372 => 0, 2373 => 0, 2374 => 0, 2375 => 0, 2376 => 0, 2377 => 0, 2378 => 0, 2379 => 0, 2380 => 0, 2381 => 0, 2382 => 0, 2383 => 0, 2384 => 0, 2385 => 0, 2386 => 0, 2387 => 0, 2388 => 0, 2389 => 0, 2390 => 0, 2391 => 0, 2392 => 0, 2393 => 0, 2394 => 0, 2395 => 0, 2396 => 0, 2397 => 0, 2398 => 0, 2399 => 0, 2400 => 0, 2401 => 1, 2402 => 1, 2403 => 1, 2404 => 1, 2405 => 1, 2406 => 1, 2407 => 1, 2408 => 1, 2409 => 1, 2410 => 1, 2411 => 1, 2412 => 0, 2413 => 0, 2414 => 0, 2415 => 0, 2416 => 0, 2417 => 0, 2418 => 0, 2419 => 0, 2420 => 0, 2421 => 0, 2422 => 0, 2423 => 0, 2424 => 0, 2425 => 0, 2426 => 0, 2427 => 0, 2428 => 0, 2429 => 0, 2430 => 0, 2431 => 0, 2432 => 0, 2433 => 0, 2434 => 0, 2435 => 0, 2436 => 0, 2437 => 0, 2438 => 0, 2439 => 0, 2440 => 0, 2441 => 0, 2442 => 0, 2443 => 0, 2444 => 0, 2445 => 0, 2446 => 0, 2447 => 0, 2448 => 0, 2449 => 0, 2450 => 0, 2451 => 0, 2452 => 0, 2453 => 0, 2454 => 0, 2455 => 0, 2456 => 0, 2457 => 0, 2458 => 0, 2459 => 1, 2460 => 1, 2461 => 1, 
2462 => 1, 2463 => 1, 2464 => 0, 2465 => 0, 2466 => 0, 2467 => 0, 2468 => 0, 2469 => 0, 2470 => 0, 2471 => 0, 2472 => 0, 2473 => 0, 2474 => 0, 2475 => 
0, 2476 => 0, 2477 => 0, 2478 => 0, 2479 => 0, 2480 => 0, 2481 => 0, 2482 => 0, 2483 => 0, 2484 => 1, 2485 => 1, 2486 => 1, 2487 => 1, 2488 => 1, 2489 
=> 0, 2490 => 0, 2491 => 0, 2492 => 0, 2493 => 0, 2494 => 0, 2495 => 0, 2496 => 0, 2497 => 0, 2498 => 0, 2499 => 0, 2500 => 0, 2501 => 0, 2502 => 0, 2503 => 0, 2504 => 1, 2505 => 1, 2506 => 1, 2507 => 1, 2508 => 1, 2509 => 1, 2510 => 1, 2511 => 1, 2512 => 1, 2513 => 1, 2514 => 1, 2515 => 1, 2516 => 0, 2517 => 0, 2518 => 0, 2519 => 0, 2520 => 0, 2521 => 0, 2522 => 0, 2523 => 0, 2524 => 0, 2525 => 0, 2526 => 0, 2527 => 0, 2528 => 0, 2529 => 0, 2530 => 0, 2531 => 0, 2532 => 0, 2533 => 0, 2534 => 0, 2535 => 0, 2536 => 1, 2537 => 1, 2538 => 1, 2539 => 1, 2540 => 1, 2541 => 1, 2542 => 1, 2543 => 1, 2544 => 1, 2545 => 1, 2546 => 1, 2547 => 0, 2548 => 0, 2549 => 0, 2550 => 0, 2551 => 0, 2552 => 0, 2553 => 0, 2554 => 0, 2555 => 1, 2556 => 1, 2557 => 1, 2558 => 1, 2559 => 1, 2560 => 1, 2561 => 1, 2562 => 1, 2563 => 1, 2564 => 1, 2565 => 1, 2566 => 1, 2567 => 0, 2568 => 0, 2569 => 0, 2570 => 0, 2571 => 0, 2572 => 0, 2573 => 0, 2574 => 0, 2575 => 0, 2576 => 0, 2577 => 0, 2578 => 0, 2579 => 0, 2580 => 0, 2581 => 0, 2582 => 0, 2583 => 0, 2584 => 0, 2585 => 0, 2586 => 0, 2587 => 0, 2588 => 0, 2589 => 0, 2590 => 0, 2591 => 0, 2592 => 0, 2593 => 0, 2594 => 0, 2595 => 0, 2596 => 0, 2597 => 0, 2598 => 0, 2599 => 0, 2600 => 0, 2601 => 1, 2602 => 1, 2603 => 1, 2604 => 1, 2605 => 1, 2606 => 1, 2607 => 1, 2608 => 1, 2609 => 1, 2610 => 1, 2611 => 1, 2612 => 0, 
2613 => 0, 2614 => 0, 2615 => 0, 2616 => 0, 2617 => 0, 2618 => 0, 2619 => 0, 2620 => 0, 2621 => 0, 2622 => 0, 2623 => 0, 2624 => 0, 2625 => 0, 2626 => 
0, 2627 => 0, 2628 => 0, 2629 => 0, 2630 => 0, 2631 => 0, 2632 => 0, 2633 => 0, 2634 => 0, 2635 => 0, 2636 => 0, 2637 => 0, 2638 => 0, 2639 => 0, 2640 
=> 0, 2641 => 0, 2642 => 0, 2643 => 0, 2644 => 0, 2645 => 0, 2646 => 0, 2647 => 0, 2648 => 0, 2649 => 0, 2650 => 0, 2651 => 0, 2652 => 1, 2653 => 1, 2654 => 1, 2655 => 1, 2656 => 1, 2657 => 1, 2658 => 1, 2659 => 1, 2660 => 1, 2661 => 1, 2662 => 1, 2663 => 1, 2664 => 0, 2665 => 0, 2666 => 0, 2667 => 0, 2668 => 0, 2669 => 0, 2670 => 0, 2671 => 0, 2672 => 0, 2673 => 0, 2674 => 0, 2675 => 0, 2676 => 0, 2677 => 0, 2678 => 0, 2679 => 0, 2680 => 0, 2681 => 0, 2682 => 0, 2683 => 0, 2684 => 1, 2685 => 1, 2686 => 1, 2687 => 1, 2688 => 1, 2689 => 1, 2690 => 1, 2691 => 1, 2692 => 1, 2693 => 1, 2694 => 1, 2695 => 1, 2696 => 0, 2697 => 0, 2698 => 0, 2699 => 0, 2700 => 0, 2701 => 0, 2702 => 0, 2703 => 0, 2704 => 1, 2705 => 1, 2706 => 1, 2707 => 1, 2708 => 1, 2709 => 1, 2710 => 1, 2711 => 1, 2712 => 1, 2713 => 1, 2714 => 1, 2715 => 1, 2716 => 1, 2717 => 1, 2718 => 1, 2719 => 1, 2720 => 1, 2721 => 1, 2722 => 0, 2723 => 0, 2724 => 0, 2725 => 0, 2726 => 0, 2727 => 0, 2728 => 0, 2729 => 0, 2730 => 1, 2731 => 1, 2732 => 1, 2733 => 1, 2734 => 1, 2735 => 1, 2736 => 1, 2737 => 1, 2738 => 1, 2739 => 1, 2740 => 1, 2741 => 1, 2742 => 1, 2743 => 1, 2744 => 1, 2745 => 1, 2746 => 1, 2747 => 0, 2748 => 0, 2749 => 0, 2750 => 0, 2751 => 0, 2752 => 0, 2753 => 0, 2754 => 0, 2755 => 1, 2756 => 1, 2757 => 1, 2758 => 1, 2759 => 1, 2760 => 1, 2761 => 1, 2762 => 1, 2763 => 1, 
2764 => 1, 2765 => 1, 2766 => 1, 2767 => 0, 2768 => 0, 2769 => 0, 2770 => 0, 2771 => 0, 2772 => 0, 2773 => 0, 2774 => 0, 2775 => 0, 2776 => 0, 2777 => 
0, 2778 => 0, 2779 => 0, 2780 => 0, 2781 => 0, 2782 => 0, 2783 => 0, 2784 => 0, 2785 => 0, 2786 => 0, 2787 => 0, 2788 => 0, 2789 => 0, 2790 => 0, 2791 
=> 0, 2792 => 0, 2793 => 0, 2794 => 0, 2795 => 0, 2796 => 0, 2797 => 0, 2798 => 0, 2799 => 0, 2800 => 0, 2801 => 1, 2802 => 1, 2803 => 1, 2804 => 1, 2805 => 1, 2806 => 1, 2807 => 1, 2808 => 1, 2809 => 1, 2810 => 1, 2811 => 1, 2812 => 0, 2813 => 0, 2814 => 0, 2815 => 0, 2816 => 0, 2817 => 0, 2818 => 0, 2819 => 0, 2820 => 0, 2821 => 0, 2822 => 0, 2823 => 0, 2824 => 0, 2825 => 0, 2826 => 0, 2827 => 0, 2828 => 0, 2829 => 0, 2830 => 0, 2831 => 0, 2832 => 0, 2833 => 0, 2834 => 0, 2835 => 0, 2836 => 0, 2837 => 0, 2838 => 0, 2839 => 0, 2840 => 0, 2841 => 0, 2842 => 0, 2843 => 0, 2844 => 0, 2845 => 0, 2846 => 0, 2847 => 0, 2848 => 0, 2849 => 0, 2850 => 0, 2851 => 0, 2852 => 1, 2853 => 1, 2854 => 1, 2855 => 1, 2856 => 1, 2857 => 1, 2858 => 1, 2859 => 1, 2860 => 1, 2861 => 1, 2862 => 1, 2863 => 1, 2864 => 0, 2865 => 0, 2866 => 0, 2867 => 0, 2868 => 0, 2869 => 0, 2870 => 0, 2871 => 0, 2872 => 0, 2873 => 0, 2874 => 0, 2875 => 0, 2876 => 0, 2877 => 0, 2878 => 0, 2879 => 0, 2880 => 0, 2881 => 0, 2882 => 0, 2883 => 0, 2884 => 1, 2885 => 1, 2886 => 1, 2887 => 1, 2888 => 1, 2889 => 1, 2890 => 1, 2891 => 1, 2892 => 1, 2893 => 1, 2894 => 1, 2895 => 1, 2896 => 0, 2897 => 0, 2898 => 0, 2899 => 0, 2900 => 0, 2901 => 0, 2902 => 0, 2903 => 0, 2904 => 1, 2905 => 1, 2906 => 1, 2907 => 1, 2908 => 1, 2909 => 1, 2910 => 1, 2911 => 1, 2912 => 1, 2913 => 1, 2914 => 1, 
2915 => 1, 2916 => 1, 2917 => 1, 2918 => 1, 2919 => 1, 2920 => 1, 2921 => 1, 2922 => 0, 2923 => 0, 2924 => 0, 2925 => 0, 2926 => 0, 2927 => 0, 2928 => 
0, 2929 => 0, 2930 => 1, 2931 => 1, 2932 => 1, 2933 => 1, 2934 => 1, 2935 => 1, 2936 => 1, 2937 => 1, 2938 => 1, 2939 => 1, 2940 => 1, 2941 => 1, 2942 
=> 1, 2943 => 1, 2944 => 1, 2945 => 1, 2946 => 1, 2947 => 0, 2948 => 0, 2949 => 0, 2950 => 0, 2951 => 0, 2952 => 0, 2953 => 0, 2954 => 0, 2955 => 1, 2956 => 1, 2957 => 1, 2958 => 1, 2959 => 1, 2960 => 1, 2961 => 1, 2962 => 1, 2963 => 1, 2964 => 1, 2965 => 1, 2966 => 1, 2967 => 0, 2968 => 0, 2969 => 0, 2970 => 0, 2971 => 0, 2972 => 0, 2973 => 0, 2974 => 0, 2975 => 0, 2976 => 0, 2977 => 0, 2978 => 0, 2979 => 0, 2980 => 0, 2981 => 0, 2982 => 0, 2983 => 0, 2984 => 0, 2985 => 0, 2986 => 0, 2987 => 0, 2988 => 0, 2989 => 0, 2990 => 0, 2991 => 0, 2992 => 0, 2993 => 0, 2994 => 0, 2995 => 0, 2996 => 0, 2997 => 0, 2998 => 0, 2999 => 0, 3000 => 0, 3001 => 1, 3002 => 1, 3003 => 1, 3004 => 1, 3005 => 1, 3006 => 1, 3007 => 1, 3008 => 1, 3009 => 1, 3010 => 1, 3011 => 1, 3012 => 0, 3013 => 0, 3014 => 0, 3015 => 0, 3016 => 0, 3017 => 0, 3018 => 0, 3019 => 0, 3020 => 0, 3021 => 0, 3022 => 0, 3023 => 0, 3024 => 0, 3025 => 0, 3026 => 0, 3027 => 0, 3028 => 0, 3029 => 0, 3030 => 0, 3031 => 0, 3032 => 0, 3033 => 0, 3034 => 0, 3035 => 0, 3036 => 0, 3037 => 0, 3038 => 0, 3039 => 0, 3040 => 0, 3041 => 0, 3042 => 0, 3043 => 0, 3044 => 0, 3045 => 0, 3046 => 0, 3047 => 0, 3048 => 0, 3049 => 0, 3050 => 0, 3051 => 0, 3052 => 1, 3053 => 1, 3054 => 1, 3055 => 1, 3056 => 1, 3057 => 1, 3058 => 1, 3059 => 1, 3060 => 1, 3061 => 1, 3062 => 1, 3063 => 1, 3064 => 0, 3065 => 0, 
3066 => 0, 3067 => 0, 3068 => 0, 3069 => 0, 3070 => 0, 3071 => 0, 3072 => 0, 3073 => 0, 3074 => 0, 3075 => 0, 3076 => 0, 3077 => 0, 3078 => 0, 3079 => 
0, 3080 => 0, 3081 => 0, 3082 => 0, 3083 => 0, 3084 => 1, 3085 => 1, 3086 => 1, 3087 => 1, 3088 => 1, 3089 => 1, 3090 => 1, 3091 => 1, 3092 => 1, 3093 
=> 1, 3094 => 1, 3095 => 1, 3096 => 0, 3097 => 0, 3098 => 0, 3099 => 0, 3100 => 0, 3101 => 0, 3102 => 0, 3103 => 0, 3104 => 1, 3105 => 1, 3106 => 1, 3107 => 1, 3108 => 1, 3109 => 1, 3110 => 1, 3111 => 1, 3112 => 1, 3113 => 1, 3114 => 1, 3115 => 1, 3116 => 1, 3117 => 1, 3118 => 1, 3119 => 1, 3120 => 1, 3121 => 1, 3122 => 0, 3123 => 0, 3124 => 0, 3125 => 0, 3126 => 0, 3127 => 0, 3128 => 0, 3129 => 0, 3130 => 1, 3131 => 1, 3132 => 1, 3133 => 1, 3134 => 1, 3135 => 1, 3136 => 1, 3137 => 1, 3138 => 1, 3139 => 1, 3140 => 1, 3141 => 1, 3142 => 1, 3143 => 1, 3144 => 1, 3145 => 1, 3146 => 1, 3147 => 0, 3148 => 0, 3149 => 0, 3150 => 0, 3151 => 0, 3152 => 0, 3153 => 0, 3154 => 0, 3155 => 1, 3156 => 1, 3157 => 1, 3158 => 1, 3159 => 1, 3160 => 1, 3161 => 1, 3162 => 1, 3163 => 1, 3164 => 1, 3165 => 1, 3166 => 1, 3167 => 0, 3168 => 0, 3169 => 0, 3170 => 0, 3171 => 0, 3172 => 0, 3173 => 0, 3174 => 0, 3175 => 0, 3176 => 0, 3177 => 0, 3178 => 0, 3179 => 0, 3180 => 0, 3181 => 0, 3182 => 0, 3183 => 0, 3184 => 0, 3185 => 0, 3186 => 0, 3187 => 0, 3188 => 0, 3189 => 0, 3190 => 0, 3191 => 0, 3192 => 0, 3193 => 0, 3194 => 0, 3195 => 0, 3196 => 0, 3197 => 0, 3198 => 0, 3199 => 0, 3200 => 0, 3201 => 1, 3202 => 1, 3203 => 1, 3204 => 1, 3205 => 1, 3206 => 1, 3207 => 1, 3208 => 1, 3209 => 1, 3210 => 1, 3211 => 1, 3212 => 0, 3213 => 0, 3214 => 0, 3215 => 0, 3216 => 0, 
3217 => 0, 3218 => 0, 3219 => 0, 3220 => 0, 3221 => 0, 3222 => 0, 3223 => 0, 3224 => 0, 3225 => 0, 3226 => 0, 3227 => 0, 3228 => 0, 3229 => 0, 3230 => 
0, 3231 => 0, 3232 => 0, 3233 => 0, 3234 => 0, 3235 => 0, 3236 => 0, 3237 => 0, 3238 => 0, 3239 => 0, 3240 => 0, 3241 => 0, 3242 => 0, 3243 => 0, 3244 
=> 0, 3245 => 0, 3246 => 0, 3247 => 0, 3248 => 0, 3249 => 0, 3250 => 0, 3251 => 0, 3252 => 1, 3253 => 1, 3254 => 1, 3255 => 1, 3256 => 1, 3257 => 1, 3258 => 1, 3259 => 1, 3260 => 1, 3261 => 1, 3262 => 1, 3263 => 1, 3264 => 0, 3265 => 0, 3266 => 0, 3267 => 0, 3268 => 0, 3269 => 0, 3270 => 0, 3271 => 0, 3272 => 0, 3273 => 0, 3274 => 0, 3275 => 0, 3276 => 0, 3277 => 0, 3278 => 0, 3279 => 0, 3280 => 0, 3281 => 0, 3282 => 0, 3283 => 0, 3284 => 1, 3285 => 1, 3286 => 1, 3287 => 1, 3288 => 1, 3289 => 1, 3290 => 1, 3291 => 1, 3292 => 1, 3293 => 1, 3294 => 1, 3295 => 1, 3296 => 0, 3297 => 0, 3298 => 0, 3299 => 0, 3300 => 0, 3301 => 0, 3302 => 0, 3303 => 0, 3304 => 1, 3305 => 1, 3306 => 1, 3307 => 1, 3308 => 1, 3309 => 1, 3310 => 1, 3311 => 1, 3312 => 1, 3313 => 1, 3314 => 1, 3315 => 1, 3316 => 1, 3317 => 1, 3318 => 1, 3319 => 1, 3320 => 1, 3321 => 1, 3322 => 0, 3323 => 0, 3324 => 0, 3325 => 0, 3326 => 0, 3327 => 0, 3328 => 0, 3329 => 0, 3330 => 1, 3331 => 1, 3332 => 1, 3333 => 1, 3334 => 1, 3335 => 1, 3336 => 1, 3337 => 1, 3338 => 1, 3339 => 1, 3340 => 1, 3341 => 1, 3342 => 1, 3343 => 1, 3344 => 1, 3345 => 1, 3346 => 1, 3347 => 0, 3348 => 0, 3349 => 0, 3350 => 0, 3351 => 0, 3352 => 0, 3353 => 0, 3354 => 0, 3355 => 1, 3356 => 1, 3357 => 1, 3358 => 1, 3359 => 1, 3360 => 1, 3361 => 1, 3362 => 1, 3363 => 1, 3364 => 1, 3365 => 1, 3366 => 1, 3367 => 0, 
3368 => 0, 3369 => 0, 3370 => 0, 3371 => 0, 3372 => 0, 3373 => 0, 3374 => 0, 3375 => 0, 3376 => 0, 3377 => 0, 3378 => 0, 3379 => 0, 3380 => 0, 3381 => 
0, 3382 => 0, 3383 => 0, 3384 => 0, 3385 => 0, 3386 => 0, 3387 => 0, 3388 => 0, 3389 => 0, 3390 => 0, 3391 => 0, 3392 => 0, 3393 => 0, 3394 => 0, 3395 
=> 0, 3396 => 0, 3397 => 0, 3398 => 0, 3399 => 0, 3400 => 0, 3401 => 1, 3402 => 1, 3403 => 1, 3404 => 1, 3405 => 1, 3406 => 1, 3407 => 1, 3408 => 1, 3409 => 1, 3410 => 1, 3411 => 1, 3412 => 0, 3413 => 0, 3414 => 0, 3415 => 0, 3416 => 0, 3417 => 0, 3418 => 0, 3419 => 0, 3420 => 0, 3421 => 0, 3422 => 0, 3423 => 0, 3424 => 0, 3425 => 0, 3426 => 0, 3427 => 0, 3428 => 0, 3429 => 0, 3430 => 0, 3431 => 0, 3432 => 0, 3433 => 0, 3434 => 0, 3435 => 0, 3436 => 0, 3437 => 0, 3438 => 0, 3439 => 0, 3440 => 0, 3441 => 0, 3442 => 0, 3443 => 0, 3444 => 0, 3445 => 0, 3446 => 0, 3447 => 0, 3448 => 0, 3449 => 0, 3450 => 0, 3451 => 0, 3452 => 1, 3453 => 1, 3454 => 1, 3455 => 1, 3456 => 1, 3457 => 1, 3458 => 1, 3459 => 1, 3460 => 1, 3461 => 1, 3462 => 1, 3463 => 1, 3464 => 0, 3465 => 0, 3466 => 0, 3467 => 0, 3468 => 0, 3469 => 0, 3470 => 0, 3471 => 0, 3472 => 0, 3473 => 0, 3474 => 0, 3475 => 0, 3476 => 0, 3477 => 0, 3478 => 0, 3479 => 0, 3480 => 0, 3481 => 0, 3482 => 0, 3483 => 0, 3484 => 1, 3485 => 1, 3486 => 1, 3487 => 1, 3488 => 1, 3489 => 1, 3490 => 1, 3491 => 1, 3492 => 1, 3493 => 1, 3494 => 1, 3495 => 1, 3496 => 0, 3497 => 0, 3498 => 0, 3499 => 0, 3500 => 0, 3501 => 0, 3502 => 0, 3503 => 0, 3504 => 1, 3505 => 1, 3506 => 1, 3507 => 1, 3508 => 1, 3509 => 1, 3510 => 1, 3511 => 1, 3512 => 1, 3513 => 1, 3514 => 1, 3515 => 1, 3516 => 1, 3517 => 1, 3518 => 1, 
3519 => 1, 3520 => 1, 3521 => 1, 3522 => 0, 3523 => 0, 3524 => 0, 3525 => 0, 3526 => 0, 3527 => 0, 3528 => 0, 3529 => 0, 3530 => 1, 3531 => 1, 3532 => 
1, 3533 => 1, 3534 => 1, 3535 => 1, 3536 => 1, 3537 => 1, 3538 => 1, 3539 => 1, 3540 => 1, 3541 => 1, 3542 => 1, 3543 => 1, 3544 => 1, 3545 => 1, 3546 
=> 1, 3547 => 0, 3548 => 0, 3549 => 0, 3550 => 0, 3551 => 0, 3552 => 0, 3553 => 0, 3554 => 0, 3555 => 1, 3556 => 1, 3557 => 1, 3558 => 1, 3559 => 1, 3560 => 1, 3561 => 1, 3562 => 1, 3563 => 1, 3564 => 1, 3565 => 1, 3566 => 1, 3567 => 0, 3568 => 0, 3569 => 0, 3570 => 0, 3571 => 0, 3572 => 0, 3573 => 0, 3574 => 0, 3575 => 0, 3576 => 0, 3577 => 0, 3578 => 0, 3579 => 0, 3580 => 0, 3581 => 0, 3582 => 0, 3583 => 0, 3584 => 0, 3585 => 0, 3586 => 0, 3587 => 0, 3588 => 0, 3589 => 0, 3590 => 0, 3591 => 0, 3592 => 0, 3593 => 0, 3594 => 0, 3595 => 0, 3596 => 0, 3597 => 0, 3598 => 0, 3599 => 0, 3600 => 0, 3601 => 1, 3602 => 1, 3603 => 1, 3604 => 1, 3605 => 1, 3606 => 1, 3607 => 1, 3608 => 1, 3609 => 1, 3610 => 1, 3611 => 1, 3612 => 0, 3613 => 0, 3614 => 0, 3615 => 0, 3616 => 0, 3617 => 0, 3618 => 0, 3619 => 0, 3620 => 0, 3621 => 0, 3622 => 0, 3623 => 0, 3624 => 0, 3625 => 0, 3626 => 0, 3627 => 0, 3628 => 0, 3629 => 0, 3630 => 0, 3631 => 0, 3632 => 0, 3633 => 0, 3634 => 0, 3635 => 0, 3636 => 0, 3637 => 0, 3638 => 0, 3639 => 0, 3640 => 0, 3641 => 0, 3642 => 0, 3643 => 0, 3644 => 0, 3645 => 0, 3646 => 0, 3647 => 0, 3648 => 0, 3649 => 0, 3650 => 0, 3651 => 0, 3652 => 1, 3653 => 1, 3654 => 1, 3655 => 1, 3656 => 1, 3657 => 1, 3658 => 1, 3659 => 1, 3660 => 1, 3661 => 1, 3662 => 1, 3663 => 1, 3664 => 0, 3665 => 0, 3666 => 0, 3667 => 0, 3668 => 0, 3669 => 0, 
3670 => 0, 3671 => 0, 3672 => 0, 3673 => 0, 3674 => 0, 3675 => 0, 3676 => 0, 3677 => 0, 3678 => 0, 3679 => 0, 3680 => 0, 3681 => 0, 3682 => 0, 3683 => 
0, 3684 => 1, 3685 => 1, 3686 => 1, 3687 => 1, 3688 => 1, 3689 => 1, 3690 => 1, 3691 => 1, 3692 => 1, 3693 => 1, 3694 => 1, 3695 => 1, 3696 => 0, 3697 
=> 0, 3698 => 0, 3699 => 0, 3700 => 0, 3701 => 0, 3702 => 0, 3703 => 0, 3704 => 1, 3705 => 1, 3706 => 1, 3707 => 1, 3708 => 1, 3709 => 1, 3710 => 1, 3711 => 1, 3712 => 1, 3713 => 1, 3714 => 1, 3715 => 1, 3716 => 1, 3717 => 1, 3718 => 1, 3719 => 1, 3720 => 1, 3721 => 1, 3722 => 0, 3723 => 0, 3724 => 0, 3725 => 0, 3726 => 0, 3727 => 0, 3728 => 0, 3729 => 0, 3730 => 1, 3731 => 1, 3732 => 1, 3733 => 1, 3734 => 1, 3735 => 1, 3736 => 1, 3737 => 1, 3738 => 1, 3739 => 1, 3740 => 1, 3741 => 1, 3742 => 1, 3743 => 1, 3744 => 1, 3745 => 1, 3746 => 1, 3747 => 0, 3748 => 0, 3749 => 0, 3750 => 0, 3751 => 0, 3752 => 0, 3753 => 0, 3754 => 0, 3755 => 1, 3756 => 1, 3757 => 1, 3758 => 1, 3759 => 1, 3760 => 1, 3761 => 1, 3762 => 1, 3763 => 1, 3764 => 1, 3765 => 1, 3766 => 1, 3767 => 0, 3768 => 0, 3769 => 0, 3770 => 0, 3771 => 0, 3772 => 0, 3773 => 0, 3774 => 0, 3775 => 0, 3776 => 0, 3777 => 0, 3778 => 0, 3779 => 0, 3780 => 0, 3781 => 0, 3782 => 0, 3783 => 0, 3784 => 0, 3785 => 0, 3786 => 0, 3787 => 0, 3788 => 0, 3789 => 0, 3790 => 0, 3791 => 0, 3792 => 0, 3793 => 0, 3794 => 0, 3795 => 0, 3796 => 0, 3797 => 0, 3798 => 0, 3799 => 0, 3800 => 0, 3801 => 1, 3802 => 1, 3803 => 1, 3804 => 1, 3805 => 1, 3806 => 1, 3807 => 1, 3808 => 1, 3809 => 1, 3810 => 1, 3811 => 1, 3812 => 0, 3813 => 0, 3814 => 0, 3815 => 0, 3816 => 0, 3817 => 0, 3818 => 0, 3819 => 0, 3820 => 0, 
3821 => 0, 3822 => 0, 3823 => 0, 3824 => 0, 3825 => 0, 3826 => 0, 3827 => 0, 3828 => 0, 3829 => 0, 3830 => 0, 3831 => 0, 3832 => 0, 3833 => 0, 3834 => 
0, 3835 => 0, 3836 => 0, 3837 => 0, 3838 => 0, 3839 => 0, 3840 => 0, 3841 => 0, 3842 => 0, 3843 => 0, 3844 => 0, 3845 => 0, 3846 => 0, 3847 => 0, 3848 
=> 0, 3849 => 0, 3850 => 0, 3851 => 0, 3852 => 1, 3853 => 1, 3854 => 1, 3855 => 1, 3856 => 1, 3857 => 1, 3858 => 1, 3859 => 1, 3860 => 1, 3861 => 1, 3862 => 1, 3863 => 1, 3864 => 0, 3865 => 0, 3866 => 0, 3867 => 0, 3868 => 0, 3869 => 0, 3870 => 0, 3871 => 0, 3872 => 0, 3873 => 0, 3874 => 0, 3875 => 0, 3876 => 0, 3877 => 0, 3878 => 0, 3879 => 0, 3880 => 0, 3881 => 0, 3882 => 0, 3883 => 0, 3884 => 1, 3885 => 1, 3886 => 1, 3887 => 1, 3888 => 1, 3889 => 1, 3890 => 1, 3891 => 1, 3892 => 1, 3893 => 1, 3894 => 1, 3895 => 1, 3896 => 0, 3897 => 0, 3898 => 0, 3899 => 0, 3900 => 0, 3901 => 0, 3902 => 0, 3903 => 0, 3904 => 1, 3905 => 1, 3906 => 1, 3907 => 1, 3908 => 1, 3909 => 1, 3910 => 1, 3911 => 1, 3912 => 1, 3913 => 1, 3914 => 1, 3915 => 1, 3916 => 0, 3917 => 0, 3918 => 0, 3919 => 0, 3920 => 0, 3921 => 0, 3922 => 0, 3923 => 0, 3924 => 0, 3925 => 0, 3926 => 0, 3927 => 0, 3928 => 0, 3929 => 0, 3930 => 0, 3931 => 0, 3932 => 0, 3933 => 0, 3934 => 0, 3935 => 0, 3936 => 1, 3937 => 1, 3938 => 1, 3939 => 1, 3940 => 1, 3941 => 1, 3942 => 1, 3943 => 1, 3944 => 1, 3945 => 1, 3946 => 1, 3947 => 0, 3948 => 0, 3949 => 0, 3950 => 0, 3951 => 0, 3952 => 0, 3953 => 0, 3954 => 0, 3955 => 1, 3956 => 1, 3957 => 1, 3958 => 1, 3959 => 1, 3960 => 1, 3961 => 1, 3962 => 1, 3963 => 1, 3964 => 1, 3965 => 1, 3966 => 1, 3967 => 0, 3968 => 0, 3969 => 0, 3970 => 0, 3971 => 0, 
3972 => 0, 3973 => 0, 3974 => 0, 3975 => 0, 3976 => 0, 3977 => 0, 3978 => 0, 3979 => 0, 3980 => 0, 3981 => 0, 3982 => 0, 3983 => 0, 3984 => 0, 3985 => 
0, 3986 => 0, 3987 => 0, 3988 => 0, 3989 => 0, 3990 => 0, 3991 => 0, 3992 => 0, 3993 => 0, 3994 => 0, 3995 => 0, 3996 => 0, 3997 => 0, 3998 => 0, 3999 
=> 0, 4000 => 0, 4001 => 1, 4002 => 1, 4003 => 1, 4004 => 1, 4005 => 1, 4006 => 1, 4007 => 1, 4008 => 1, 4009 => 1, 4010 => 1, 4011 => 1, 4012 => 0, 4013 => 0, 4014 => 0, 4015 => 0, 4016 => 0, 4017 => 0, 4018 => 0, 4019 => 0, 4020 => 1, 4021 => 1, 4022 => 1, 4023 => 1, 4024 => 1, 4025 => 1, 4026 => 1, 4027 => 1, 4028 => 1, 4029 => 1, 4030 => 1, 4031 => 1, 4032 => 1, 4033 => 1, 4034 => 1, 4035 => 1, 4036 => 1, 4037 => 1, 4038 => 1, 4039 => 1, 4040 => 1, 4041 => 1, 4042 => 1, 4043 => 1, 4044 => 0, 4045 => 0, 4046 => 0, 4047 => 0, 4048 => 0, 4049 => 0, 4050 => 0, 4051 => 0, 4052 => 1, 4053 => 1, 4054 => 1, 4055 => 1, 4056 => 1, 4057 => 1, 4058 => 1, 4059 => 1, 4060 => 1, 4061 => 1, 4062 => 1, 4063 => 1, 4064 => 0, 4065 => 0, 4066 => 0, 4067 => 0, 4068 => 0, 4069 => 0, 4070 => 0, 4071 => 0, 4072 => 0, 4073 => 0, 4074 => 0, 4075 => 0, 4076 => 0, 4077 => 0, 4078 => 0, 4079 => 0, 4080 => 0, 4081 => 0, 4082 => 0, 4083 => 0, 4084 => 1, 4085 => 1, 4086 => 1, 4087 => 1, 4088 => 1, 4089 => 1, 4090 => 1, 4091 => 1, 4092 => 1, 4093 => 1, 4094 => 1, 4095 => 1, 4096 => 0, 4097 => 0, 4098 => 0, 4099 => 0, 4100 => 0, 4101 => 0, 4102 => 0, 4103 => 0, 4104 => 1, 4105 => 1, 4106 => 1, 4107 => 1, 4108 => 1, 4109 => 1, 4110 => 1, 4111 => 1, 4112 => 1, 4113 => 1, 4114 => 1, 4115 => 1, 4116 => 0, 4117 => 0, 4118 => 0, 4119 => 0, 4120 => 0, 4121 => 0, 4122 => 0, 
4123 => 1, 4124 => 1, 4125 => 1, 4126 => 1, 4127 => 1, 4128 => 0, 4129 => 0, 4130 => 0, 4131 => 0, 4132 => 0, 4133 => 0, 4134 => 0, 4135 => 0, 4136 => 
1, 4137 => 1, 4138 => 1, 4139 => 1, 4140 => 1, 4141 => 1, 4142 => 1, 4143 => 1, 4144 => 1, 4145 => 1, 4146 => 1, 4147 => 0, 4148 => 0, 4149 => 0, 4150 
=> 0, 4151 => 0, 4152 => 0, 4153 => 0, 4154 => 0, 4155 => 1, 4156 => 1, 4157 => 1, 4158 => 1, 4159 => 1, 4160 => 1, 4161 => 1, 4162 => 1, 4163 => 1, 4164 => 1, 4165 => 1, 4166 => 1, 4167 => 1, 4168 => 1, 4169 => 1, 4170 => 1, 4171 => 1, 4172 => 1, 4173 => 1, 4174 => 1, 4175 => 1, 4176 => 1, 4177 => 1, 4178 => 1, 4179 => 1, 4180 => 1, 4181 => 1, 4182 => 1, 4183 => 1, 4184 => 1, 4185 => 1, 4186 => 1, 4187 => 1, 4188 => 1, 4189 => 1, 4190 => 1, 4191 => 1, 4192 => 1, 4193 => 0, 4194 => 0, 4195 => 0, 4196 => 0, 4197 => 0, 4198 => 0, 4199 => 0, 4200 => 0, 4201 => 1, 4202 => 1, 4203 => 1, 4204 => 1, 4205 => 1, 4206 => 1, 4207 => 1, 4208 => 1, 4209 => 1, 4210 => 1, 4211 => 1, 4212 => 0, 4213 => 0, 4214 => 0, 4215 => 0, 4216 => 0, 4217 => 0, 4218 => 0, 4219 => 0, 4220 => 1, 4221 => 1, 4222 => 1, 4223 => 1, 4224 => 1, 4225 => 1, 4226 => 1, 4227 => 1, 4228 => 1, 4229 => 1, 4230 => 1, 4231 => 1, 4232 => 1, 4233 => 1, 4234 => 1, 4235 => 1, 4236 => 1, 4237 => 1, 4238 => 1, 4239 => 1, 4240 => 1, 4241 => 1, 4242 => 1, 4243 => 1, 4244 => 0, 4245 => 0, 4246 => 0, 4247 => 0, 4248 => 0, 4249 => 0, 4250 => 0, 4251 => 0, 4252 => 1, 4253 => 1, 4254 => 1, 4255 => 1, 4256 => 1, 4257 => 1, 4258 => 1, 4259 => 1, 4260 => 1, 4261 => 1, 4262 => 1, 4263 => 1, 4264 => 0, 4265 => 0, 4266 => 0, 4267 => 0, 4268 => 0, 4269 => 0, 4270 => 0, 4271 => 0, 4272 => 0, 4273 => 0, 
4274 => 0, 4275 => 0, 4276 => 0, 4277 => 0, 4278 => 0, 4279 => 0, 4280 => 0, 4281 => 0, 4282 => 0, 4283 => 0, 4284 => 1, 4285 => 1, 4286 => 1, 4287 => 
1, 4288 => 1, 4289 => 1, 4290 => 1, 4291 => 1, 4292 => 1, 4293 => 1, 4294 => 1, 4295 => 1, 4296 => 0, 4297 => 0, 4298 => 0, 4299 => 0, 4300 => 0, 4301 
=> 0, 4302 => 0, 4303 => 0, 4304 => 1, 4305 => 1, 4306 => 1, 4307 => 1, 4308 => 1, 4309 => 1, 4310 => 1, 4311 => 1, 4312 => 1, 4313 => 1, 4314 => 1, 4315 => 1, 4316 => 0, 4317 => 0, 4318 => 0, 4319 => 0, 4320 => 0, 4321 => 0, 4322 => 0, 4323 => 1, 4324 => 1, 4325 => 1, 4326 => 1, 4327 => 1, 4328 => 0, 4329 => 0, 4330 => 0, 4331 => 0, 4332 => 0, 4333 => 0, 4334 => 0, 4335 => 0, 4336 => 1, 4337 => 1, 4338 => 1, 4339 => 1, 4340 => 1, 4341 => 1, 4342 => 1, 4343 => 1, 4344 => 1, 4345 => 1, 4346 => 1, 4347 => 0, 4348 => 0, 4349 => 0, 4350 => 0, 4351 => 0, 4352 => 0, 4353 => 0, 4354 => 0, 4355 => 1, 4356 => 1, 4357 => 1, 4358 => 1, 4359 => 1, 4360 => 1, 4361 => 1, 4362 => 1, 4363 => 1, 4364 => 1, 4365 => 1, 4366 => 1, 4367 => 1, 4368 => 1, 4369 => 1, 4370 => 1, 4371 => 1, 4372 => 1, 4373 => 1, 4374 => 1, 4375 => 1, 4376 => 1, 4377 => 1, 4378 => 1, 4379 => 1, 4380 => 1, 4381 => 1, 4382 => 1, 4383 => 1, 4384 => 1, 4385 => 1, 4386 => 1, 4387 => 1, 4388 => 1, 4389 => 1, 4390 => 1, 4391 => 1, 4392 => 1, 4393 => 0, 4394 => 0, 4395 => 0, 4396 => 0, 4397 => 0, 4398 => 0, 4399 => 0, 4400 => 0, 4401 => 1, 4402 => 1, 4403 => 1, 4404 => 1, 4405 => 1, 4406 => 1, 4407 => 1, 4408 => 1, 4409 => 1, 4410 => 1, 4411 => 1, 4412 => 0, 4413 => 0, 4414 => 0, 4415 => 0, 4416 => 0, 4417 => 0, 4418 => 0, 4419 => 0, 4420 => 1, 4421 => 1, 4422 => 1, 4423 => 1, 4424 => 1, 
4425 => 1, 4426 => 1, 4427 => 1, 4428 => 1, 4429 => 1, 4430 => 1, 4431 => 1, 4432 => 1, 4433 => 1, 4434 => 1, 4435 => 1, 4436 => 1, 4437 => 1, 4438 => 
1, 4439 => 1, 4440 => 1, 4441 => 1, 4442 => 1, 4443 => 1, 4444 => 0, 4445 => 0, 4446 => 0, 4447 => 0, 4448 => 0, 4449 => 0, 4450 => 0, 4451 => 0, 4452 
=> 1, 4453 => 1, 4454 => 1, 4455 => 1, 4456 => 1, 4457 => 1, 4458 => 1, 4459 => 1, 4460 => 1, 4461 => 1, 4462 => 1, 4463 => 1, 4464 => 0, 4465 => 0, 4466 => 0, 4467 => 0, 4468 => 0, 4469 => 0, 4470 => 0, 4471 => 0, 4472 => 0, 4473 => 0, 4474 => 0, 4475 => 0, 4476 => 0, 4477 => 0, 4478 => 0, 4479 => 0, 4480 => 0, 4481 => 0, 4482 => 0, 4483 => 0, 4484 => 1, 4485 => 1, 4486 => 1, 4487 => 1, 4488 => 1, 4489 => 1, 4490 => 1, 4491 => 1, 4492 => 1, 4493 => 1, 4494 => 1, 4495 => 1, 4496 => 0, 4497 => 0, 4498 => 0, 4499 => 0, 4500 => 0, 4501 => 0, 4502 => 0, 4503 => 0, 4504 => 1, 4505 => 1, 4506 => 1, 4507 => 1, 4508 => 1, 4509 => 1, 4510 => 1, 4511 => 1, 4512 => 1, 4513 => 1, 4514 => 1, 4515 => 1, 4516 => 0, 4517 => 0, 4518 => 0, 4519 => 0, 4520 => 0, 4521 => 0, 4522 => 0, 4523 => 1, 4524 => 1, 4525 => 1, 4526 => 1, 4527 => 1, 4528 => 0, 4529 => 0, 4530 => 0, 4531 => 0, 4532 => 0, 4533 => 0, 4534 => 0, 4535 => 0, 4536 => 1, 4537 => 1, 4538 => 1, 4539 => 1, 4540 => 1, 4541 => 1, 4542 => 1, 4543 => 1, 4544 => 1, 4545 => 1, 4546 => 1, 4547 => 0, 4548 => 0, 4549 => 0, 4550 => 0, 4551 => 0, 4552 => 0, 4553 => 0, 4554 => 0, 4555 => 1, 4556 => 1, 4557 => 1, 4558 => 1, 4559 => 1, 4560 => 1, 4561 => 1, 4562 => 1, 4563 => 1, 4564 => 1, 4565 => 1, 4566 => 1, 4567 => 1, 4568 => 1, 4569 => 1, 4570 => 1, 4571 => 1, 4572 => 1, 4573 => 1, 4574 => 1, 4575 => 1, 
4576 => 1, 4577 => 1, 4578 => 1, 4579 => 1, 4580 => 1, 4581 => 1, 4582 => 1, 4583 => 1, 4584 => 1, 4585 => 1, 4586 => 1, 4587 => 1, 4588 => 1, 4589 => 
1, 4590 => 1, 4591 => 1, 4592 => 1, 4593 => 0, 4594 => 0, 4595 => 0, 4596 => 0, 4597 => 0, 4598 => 0, 4599 => 0, 4600 => 0, 4601 => 1, 4602 => 1, 4603 
=> 1, 4604 => 1, 4605 => 1, 4606 => 1, 4607 => 1, 4608 => 1, 4609 => 1, 4610 => 1, 4611 => 1, 4612 => 0, 4613 => 0, 4614 => 0, 4615 => 0, 4616 => 0, 4617 => 0, 4618 => 0, 4619 => 0, 4620 => 1, 4621 => 1, 4622 => 1, 4623 => 1, 4624 => 1, 4625 => 1, 4626 => 1, 4627 => 1, 4628 => 1, 4629 => 1, 4630 => 1, 4631 => 1, 4632 => 1, 4633 => 1, 4634 => 1, 4635 => 1, 4636 => 1, 4637 => 1, 4638 => 1, 4639 => 1, 4640 => 1, 4641 => 1, 4642 => 1, 4643 => 1, 4644 => 0, 4645 => 0, 4646 => 0, 4647 => 0, 4648 => 0, 4649 => 0, 4650 => 0, 4651 => 0, 4652 => 1, 4653 => 1, 4654 => 1, 4655 => 1, 4656 => 1, 4657 => 1, 4658 => 1, 4659 => 1, 4660 => 1, 4661 => 1, 4662 => 1, 4663 => 1, 4664 => 0, 4665 => 0, 4666 => 0, 4667 => 0, 4668 => 0, 4669 => 0, 4670 => 0, 4671 => 0, 4672 => 0, 4673 => 0, 4674 => 0, 4675 => 0, 4676 => 0, 4677 => 0, 4678 => 0, 4679 => 0, 4680 => 0, 4681 => 0, 4682 => 0, 4683 => 0, 4684 => 1, 4685 => 1, 4686 => 1, 4687 => 1, 4688 => 1, 4689 => 1, 4690 => 1, 4691 => 1, 4692 => 1, 4693 => 1, 4694 => 1, 4695 => 1, 4696 => 0, 4697 => 0, 4698 => 0, 4699 => 0, 4700 => 0, 4701 => 0, 4702 => 0, 4703 => 0, 4704 => 1, 4705 => 1, 4706 => 1, 4707 => 1, 4708 => 1, 4709 => 1, 4710 => 1, 4711 => 1, 4712 => 1, 4713 => 1, 4714 => 1, 4715 => 1, 4716 => 0, 4717 => 0, 4718 => 0, 4719 => 0, 4720 => 0, 4721 => 0, 4722 => 0, 4723 => 1, 4724 => 1, 4725 => 1, 4726 => 1, 
4727 => 1, 4728 => 0, 4729 => 0, 4730 => 0, 4731 => 0, 4732 => 0, 4733 => 0, 4734 => 0, 4735 => 0, 4736 => 1, 4737 => 1, 4738 => 1, 4739 => 1, 4740 => 
1, 4741 => 1, 4742 => 1, 4743 => 1, 4744 => 1, 4745 => 1, 4746 => 1, 4747 => 0, 4748 => 0, 4749 => 0, 4750 => 0, 4751 => 0, 4752 => 0, 4753 => 0, 4754 
=> 0, 4755 => 1, 4756 => 1, 4757 => 1, 4758 => 1, 4759 => 1, 4760 => 1, 4761 => 1, 4762 => 1, 4763 => 1, 4764 => 1, 4765 => 1, 4766 => 1, 4767 => 1, 4768 => 1, 4769 => 1, 4770 => 1, 4771 => 1, 4772 => 1, 4773 => 1, 4774 => 1, 4775 => 1, 4776 => 1, 4777 => 1, 4778 => 1, 4779 => 1, 4780 => 1, 4781 => 1, 4782 => 1, 4783 => 1, 4784 => 1, 4785 => 1, 4786 => 1, 4787 => 1, 4788 => 1, 4789 => 1, 4790 => 1, 4791 => 1, 4792 => 1, 4793 => 0, 4794 => 0, 4795 => 0, 4796 => 0, 4797 => 0, 4798 => 0, 4799 => 0, 4800 => 0, 4801 => 1, 4802 => 1, 4803 => 1, 4804 => 1, 4805 => 1, 4806 => 1, 4807 => 1, 4808 => 1, 4809 => 1, 4810 => 1, 4811 => 1, 4812 => 0, 4813 => 0, 4814 => 0, 4815 => 0, 4816 => 0, 4817 => 0, 4818 => 0, 4819 => 0, 4820 => 1, 4821 => 1, 4822 => 1, 4823 => 1, 4824 => 1, 4825 => 1, 4826 => 1, 4827 => 1, 4828 => 1, 4829 => 1, 4830 => 1, 4831 => 1, 4832 => 1, 4833 => 1, 4834 => 1, 4835 => 1, 4836 => 1, 4837 => 1, 4838 => 1, 4839 => 1, 4840 => 1, 4841 => 1, 4842 => 1, 4843 => 1, 4844 => 0, 4845 => 0, 4846 => 0, 4847 => 0, 4848 => 0, 4849 => 0, 4850 => 0, 4851 => 0, 4852 => 1, 4853 => 1, 4854 => 1, 4855 => 1, 4856 => 1, 4857 => 1, 4858 => 1, 4859 => 1, 4860 => 1, 4861 => 1, 4862 => 1, 4863 => 1, 4864 => 0, 4865 => 0, 4866 => 0, 4867 => 0, 4868 => 0, 4869 => 0, 4870 => 0, 4871 => 0, 4872 => 0, 4873 => 0, 4874 => 0, 4875 => 0, 4876 => 0, 4877 => 0, 
4878 => 0, 4879 => 0, 4880 => 0, 4881 => 0, 4882 => 0, 4883 => 0, 4884 => 1, 4885 => 1, 4886 => 1, 4887 => 1, 4888 => 1, 4889 => 1, 4890 => 1, 4891 => 
1, 4892 => 1, 4893 => 1, 4894 => 1, 4895 => 1, 4896 => 0, 4897 => 0, 4898 => 0, 4899 => 0, 4900 => 0, 4901 => 0, 4902 => 0, 4903 => 0, 4904 => 1, 4905 
=> 1, 4906 => 1, 4907 => 1, 4908 => 1, 4909 => 1, 4910 => 1, 4911 => 1, 4912 => 1, 4913 => 1, 4914 => 1, 4915 => 1, 4916 => 0, 4917 => 0, 4918 => 0, 4919 => 0, 4920 => 0, 4921 => 0, 4922 => 0, 4923 => 1, 4924 => 1, 4925 => 1, 4926 => 1, 4927 => 1, 4928 => 0, 4929 => 0, 4930 => 0, 4931 => 0, 4932 => 0, 4933 => 0, 4934 => 0, 4935 => 0, 4936 => 1, 4937 => 1, 4938 => 1, 4939 => 1, 4940 => 1, 4941 => 1, 4942 => 1, 4943 => 1, 4944 => 1, 4945 => 1, 4946 => 1, 4947 => 0, 4948 => 0, 4949 => 0, 4950 => 0, 4951 => 0, 4952 => 0, 4953 => 0, 4954 => 0, 4955 => 1, 4956 => 1, 4957 => 1, 4958 => 1, 4959 => 1, 4960 => 1, 4961 => 1, 4962 => 1, 4963 => 1, 4964 => 1, 4965 => 1, 4966 => 1, 4967 => 1, 4968 => 1, 4969 => 1, 4970 => 1, 4971 => 1, 4972 => 1, 4973 => 1, 4974 => 1, 4975 => 1, 4976 => 1, 4977 => 1, 4978 => 1, 4979 => 1, 4980 => 1, 4981 => 1, 4982 => 1, 4983 => 1, 4984 => 1, 4985 => 1, 4986 => 1, 4987 => 1, 4988 => 1, 4989 => 1, 4990 => 1, 4991 => 1, 4992 => 1, 4993 => 0, 4994 => 0, 4995 => 0, 4996 => 0, 4997 => 0, 4998 => 0, 4999 => 0, 5000 => 0, 5001 => 1, 5002 => 1, 5003 => 1, 5004 => 1, 5005 => 1, 5006 => 1, 5007 => 1, 5008 => 1, 5009 => 1, 5010 => 1, 5011 => 1, 5012 => 0, 5013 => 0, 5014 => 0, 5015 => 0, 5016 => 0, 5017 => 0, 5018 => 0, 5019 => 0, 5020 => 0, 5021 => 0, 5022 => 0, 5023 => 0, 5024 => 0, 5025 => 0, 5026 => 0, 5027 => 0, 5028 => 0, 
5029 => 0, 5030 => 0, 5031 => 0, 5032 => 0, 5033 => 1, 5034 => 1, 5035 => 1, 5036 => 1, 5037 => 1, 5038 => 1, 5039 => 1, 5040 => 1, 5041 => 1, 5042 => 
1, 5043 => 1, 5044 => 0, 5045 => 0, 5046 => 0, 5047 => 0, 5048 => 0, 5049 => 0, 5050 => 0, 5051 => 0, 5052 => 1, 5053 => 1, 5054 => 1, 5055 => 1, 5056 
=> 1, 5057 => 1, 5058 => 1, 5059 => 1, 5060 => 1, 5061 => 1, 5062 => 1, 5063 => 1, 5064 => 0, 5065 => 0, 5066 => 0, 5067 => 0, 5068 => 0, 5069 => 0, 5070 => 0, 5071 => 0, 5072 => 0, 5073 => 0, 5074 => 0, 5075 => 0, 5076 => 0, 5077 => 0, 5078 => 0, 5079 => 0, 5080 => 0, 5081 => 0, 5082 => 0, 5083 => 0, 5084 => 1, 5085 => 1, 5086 => 1, 5087 => 1, 5088 => 1, 5089 => 1, 5090 => 1, 5091 => 1, 5092 => 1, 5093 => 1, 5094 => 1, 5095 => 1, 5096 => 0, 5097 => 0, 5098 => 0, 5099 => 0, 5100 => 0, 5101 => 0, 5102 => 0, 5103 => 0, 5104 => 1, 5105 => 1, 5106 => 1, 5107 => 1, 5108 => 1, 5109 => 1, 5110 => 1, 5111 => 1, 5112 => 1, 5113 => 1, 5114 => 1, 5115 => 1, 5116 => 0, 5117 => 0, 5118 => 0, 5119 => 0, 5120 => 0, 5121 => 0, 5122 => 0, 5123 => 0, 5124 => 0, 5125 => 0, 5126 => 0, 5127 => 0, 5128 => 0, 5129 => 0, 5130 => 0, 5131 => 0, 5132 => 0, 5133 => 0, 5134 => 0, 5135 => 0, 5136 => 1, 5137 => 1, 5138 => 1, 5139 => 1, 5140 => 1, 5141 => 1, 5142 => 1, 5143 => 1, 5144 => 1, 5145 => 1, 5146 => 1, 5147 => 0, 5148 => 0, 5149 => 0, 5150 => 0, 5151 => 0, 5152 => 0, 5153 => 0, 5154 => 0, 5155 => 1, 5156 => 1, 5157 => 1, 5158 => 1, 5159 => 1, 5160 => 1, 5161 => 1, 5162 => 1, 5163 => 1, 5164 => 1, 5165 => 1, 5166 => 1, 5167 => 0, 5168 => 0, 5169 => 0, 5170 => 0, 5171 => 0, 5172 => 0, 5173 => 0, 5174 => 0, 5175 => 0, 5176 => 0, 5177 => 0, 5178 => 0, 5179 => 0, 
5180 => 0, 5181 => 0, 5182 => 0, 5183 => 0, 5184 => 0, 5185 => 0, 5186 => 0, 5187 => 0, 5188 => 0, 5189 => 0, 5190 => 0, 5191 => 0, 5192 => 0, 5193 => 
0, 5194 => 0, 5195 => 0, 5196 => 0, 5197 => 0, 5198 => 0, 5199 => 0, 5200 => 0, 5201 => 1, 5202 => 1, 5203 => 1, 5204 => 1, 5205 => 1, 5206 => 1, 5207 
=> 1, 5208 => 1, 5209 => 1, 5210 => 1, 5211 => 1, 5212 => 0, 5213 => 0, 5214 => 0, 5215 => 0, 5216 => 0, 5217 => 0, 5218 => 0, 5219 => 0, 5220 => 0, 5221 => 0, 5222 => 0, 5223 => 0, 5224 => 0, 5225 => 0, 5226 => 0, 5227 => 0, 5228 => 0, 5229 => 0, 5230 => 0, 5231 => 0, 5232 => 0, 5233 => 1, 5234 => 1, 5235 => 1, 5236 => 1, 5237 => 1, 5238 => 1, 5239 => 1, 5240 => 1, 5241 => 1, 5242 => 1, 5243 => 1, 5244 => 0, 5245 => 0, 5246 => 0, 5247 => 0, 5248 => 0, 5249 => 0, 5250 => 0, 5251 => 0, 5252 => 1, 5253 => 1, 5254 => 1, 5255 => 1, 5256 => 1, 5257 => 1, 5258 => 1, 5259 => 1, 5260 => 1, 5261 => 1, 5262 => 1, 5263 => 1, 5264 => 1, 5265 => 1, 5266 => 1, 5267 => 1, 5268 => 1, 5269 => 1, 5270 => 1, 5271 => 1, 5272 => 1, 5273 => 1, 5274 => 1, 5275 => 1, 5276 => 1, 5277 => 1, 5278 => 1, 5279 => 1, 5280 => 1, 5281 => 1, 5282 => 1, 5283 => 1, 5284 => 1, 5285 => 1, 5286 => 1, 5287 => 1, 5288 => 1, 5289 => 1, 5290 => 1, 5291 => 1, 5292 => 1, 5293 => 1, 5294 => 1, 5295 => 1, 5296 => 0, 5297 => 0, 5298 => 0, 5299 => 0, 5300 => 0, 5301 => 0, 5302 => 0, 5303 => 0, 5304 => 1, 5305 => 1, 5306 => 1, 5307 => 1, 5308 => 1, 5309 => 1, 5310 => 1, 5311 => 1, 5312 => 1, 5313 => 1, 5314 => 1, 5315 => 1, 5316 => 0, 5317 => 0, 5318 => 0, 5319 => 0, 5320 => 0, 5321 => 0, 5322 => 0, 5323 => 0, 5324 => 0, 5325 => 0, 5326 => 0, 5327 => 0, 5328 => 0, 5329 => 0, 5330 => 0, 
5331 => 0, 5332 => 0, 5333 => 0, 5334 => 0, 5335 => 0, 5336 => 1, 5337 => 1, 5338 => 1, 5339 => 1, 5340 => 1, 5341 => 1, 5342 => 1, 5343 => 1, 5344 => 
1, 5345 => 1, 5346 => 1, 5347 => 0, 5348 => 0, 5349 => 0, 5350 => 0, 5351 => 0, 5352 => 0, 5353 => 0, 5354 => 0, 5355 => 1, 5356 => 1, 5357 => 1, 5358 
=> 1, 5359 => 1, 5360 => 1, 5361 => 1, 5362 => 1, 5363 => 1, 5364 => 1, 5365 => 1, 5366 => 1, 5367 => 0, 5368 => 0, 5369 => 0, 5370 => 0, 5371 => 0, 5372 => 0, 5373 => 0, 5374 => 0, 5375 => 0, 5376 => 0, 5377 => 0, 5378 => 0, 5379 => 0, 5380 => 0, 5381 => 0, 5382 => 0, 5383 => 0, 5384 => 0, 5385 => 0, 5386 => 0, 5387 => 0, 5388 => 0, 5389 => 0, 5390 => 0, 5391 => 0, 5392 => 0, 5393 => 0, 5394 => 0, 5395 => 0, 5396 => 0, 5397 => 0, 5398 => 0, 5399 => 0, 5400 => 0, 5401 => 1, 5402 => 1, 5403 => 1, 5404 => 1, 5405 => 1, 5406 => 1, 5407 => 1, 5408 => 1, 5409 => 1, 5410 => 1, 5411 => 1, 5412 => 0, 5413 => 0, 5414 => 0, 5415 => 0, 5416 => 0, 5417 => 0, 5418 => 0, 5419 => 0, 5420 => 0, 5421 => 0, 5422 => 0, 5423 => 0, 5424 => 0, 5425 => 0, 5426 => 0, 5427 => 0, 5428 => 0, 5429 => 0, 5430 => 0, 5431 => 0, 5432 => 0, 5433 => 1, 5434 => 1, 5435 => 1, 5436 => 1, 5437 => 1, 5438 => 1, 5439 => 1, 5440 => 1, 5441 => 1, 5442 => 1, 5443 => 1, 5444 => 0, 5445 => 0, 5446 => 0, 5447 => 0, 5448 => 0, 5449 => 0, 5450 => 0, 5451 => 0, 5452 => 1, 5453 => 1, 5454 => 1, 5455 => 1, 5456 => 1, 5457 => 1, 5458 => 1, 5459 => 1, 5460 => 1, 5461 => 1, 5462 => 1, 5463 => 1, 5464 => 1, 5465 => 1, 5466 => 1, 5467 => 1, 5468 => 1, 5469 => 1, 5470 => 1, 5471 => 1, 5472 => 1, 5473 => 1, 5474 => 1, 5475 => 1, 5476 => 1, 5477 => 1, 5478 => 1, 5479 => 1, 5480 => 1, 5481 => 1, 
5482 => 1, 5483 => 1, 5484 => 1, 5485 => 1, 5486 => 1, 5487 => 1, 5488 => 1, 5489 => 1, 5490 => 1, 5491 => 1, 5492 => 1, 5493 => 1, 5494 => 1, 5495 => 
1, 5496 => 0, 5497 => 0, 5498 => 0, 5499 => 0, 5500 => 0, 5501 => 0, 5502 => 0, 5503 => 0, 5504 => 1, 5505 => 1, 5506 => 1, 5507 => 1, 5508 => 1, 5509 
=> 1, 5510 => 1, 5511 => 1, 5512 => 1, 5513 => 1, 5514 => 1, 5515 => 1, 5516 => 0, 5517 => 0, 5518 => 0, 5519 => 0, 5520 => 0, 5521 => 0, 5522 => 0, 5523 => 0, 5524 => 0, 5525 => 0, 5526 => 0, 5527 => 0, 5528 => 0, 5529 => 0, 5530 => 0, 5531 => 0, 5532 => 0, 5533 => 0, 5534 => 0, 5535 => 0, 5536 => 1, 5537 => 1, 5538 => 1, 5539 => 1, 5540 => 1, 5541 => 1, 5542 => 1, 5543 => 1, 5544 => 1, 5545 => 1, 5546 => 1, 5547 => 0, 5548 => 0, 5549 => 0, 5550 => 0, 5551 => 0, 5552 => 0, 5553 => 0, 5554 => 0, 5555 => 1, 5556 => 1, 5557 => 1, 5558 => 1, 5559 => 1, 5560 => 1, 5561 => 1, 5562 => 1, 5563 => 1, 5564 => 1, 5565 => 1, 5566 => 1, 5567 => 0, 5568 => 0, 5569 => 0, 5570 => 0, 5571 => 0, 5572 => 0, 5573 => 0, 5574 => 0, 5575 => 0, 5576 => 0, 5577 => 0, 5578 => 0, 5579 => 0, 5580 => 0, 5581 => 0, 5582 => 0, 5583 => 0, 5584 => 0, 5585 => 0, 5586 => 0, 5587 => 0, 5588 => 0, 5589 => 0, 5590 => 0, 5591 => 0, 5592 => 0, 5593 => 0, 5594 => 0, 5595 => 0, 5596 => 0, 5597 => 0, 5598 => 0, 5599 => 0, 5600 => 0, 5601 => 1, 5602 => 1, 5603 => 1, 5604 => 1, 5605 => 1, 5606 => 1, 5607 => 1, 5608 => 1, 5609 => 1, 5610 => 1, 5611 => 1, 5612 => 0, 5613 => 0, 5614 => 0, 5615 => 0, 5616 => 0, 5617 => 0, 5618 => 0, 5619 => 0, 5620 => 0, 5621 => 0, 5622 => 0, 5623 => 0, 5624 => 0, 5625 => 0, 5626 => 0, 5627 => 0, 5628 => 0, 5629 => 0, 5630 => 0, 5631 => 0, 5632 => 0, 
5633 => 1, 5634 => 1, 5635 => 1, 5636 => 1, 5637 => 1, 5638 => 1, 5639 => 1, 5640 => 1, 5641 => 1, 5642 => 1, 5643 => 1, 5644 => 0, 5645 => 0, 5646 => 
0, 5647 => 0, 5648 => 0, 5649 => 0, 5650 => 0, 5651 => 0, 5652 => 1, 5653 => 1, 5654 => 1, 5655 => 1, 5656 => 1, 5657 => 1, 5658 => 1, 5659 => 1, 5660 
=> 1, 5661 => 1, 5662 => 1, 5663 => 1, 5664 => 1, 5665 => 1, 5666 => 1, 5667 => 1, 5668 => 1, 5669 => 1, 5670 => 1, 5671 => 1, 5672 => 1, 5673 => 1, 5674 => 1, 5675 => 1, 5676 => 1, 5677 => 1, 5678 => 1, 5679 => 1, 5680 => 1, 5681 => 1, 5682 => 1, 5683 => 1, 5684 => 1, 5685 => 1, 5686 => 1, 5687 => 1, 5688 => 1, 5689 => 1, 5690 => 1, 5691 => 1, 5692 => 1, 5693 => 1, 5694 => 1, 5695 => 1, 5696 => 0, 5697 => 0, 5698 => 0, 5699 => 0, 5700 => 0, 5701 => 0, 5702 => 0, 5703 => 0, 5704 => 1, 5705 => 1, 5706 => 1, 5707 => 1, 5708 => 1, 5709 => 1, 5710 => 1, 5711 => 1, 5712 => 1, 5713 => 1, 5714 => 1, 5715 => 1, 5716 => 0, 5717 => 0, 5718 => 0, 5719 => 0, 5720 => 0, 5721 => 0, 5722 => 0, 5723 => 0, 5724 => 0, 5725 => 0, 5726 => 0, 5727 => 0, 5728 => 0, 5729 => 0, 5730 => 0, 5731 => 0, 5732 => 0, 5733 => 0, 5734 => 0, 5735 => 0, 5736 => 1, 5737 => 1, 5738 => 1, 5739 => 1, 5740 => 1, 5741 => 1, 5742 => 1, 5743 => 1, 5744 => 1, 5745 => 1, 5746 => 1, 5747 => 0, 5748 => 0, 5749 => 0, 5750 => 0, 5751 => 0, 5752 => 0, 5753 => 0, 5754 => 0, 5755 => 1, 5756 => 1, 5757 => 1, 5758 => 1, 5759 => 1, 5760 => 1, 5761 => 1, 5762 => 1, 5763 => 1, 5764 => 1, 5765 => 1, 5766 => 1, 5767 => 0, 5768 => 0, 5769 => 0, 5770 => 0, 5771 => 0, 5772 => 0, 5773 => 0, 5774 => 0, 5775 => 0, 5776 => 0, 5777 => 0, 5778 => 0, 5779 => 0, 5780 => 0, 5781 => 0, 5782 => 0, 5783 => 0, 
5784 => 0, 5785 => 0, 5786 => 0, 5787 => 0, 5788 => 0, 5789 => 0, 5790 => 0, 5791 => 0, 5792 => 0, 5793 => 0, 5794 => 0, 5795 => 0, 5796 => 0, 5797 => 
0, 5798 => 0, 5799 => 0, 5800 => 0, 5801 => 1, 5802 => 1, 5803 => 1, 5804 => 1, 5805 => 1, 5806 => 1, 5807 => 1, 5808 => 1, 5809 => 1, 5810 => 1, 5811 
=> 1, 5812 => 0, 5813 => 0, 5814 => 0, 5815 => 0, 5816 => 0, 5817 => 0, 5818 => 0, 5819 => 0, 5820 => 0, 5821 => 0, 5822 => 0, 5823 => 0, 5824 => 0, 5825 => 0, 5826 => 0, 5827 => 0, 5828 => 0, 5829 => 0, 5830 => 0, 5831 => 0, 5832 => 0, 5833 => 1, 5834 => 1, 5835 => 1, 5836 => 1, 5837 => 1, 5838 => 1, 5839 => 1, 5840 => 1, 5841 => 1, 5842 => 1, 5843 => 1, 5844 => 0, 5845 => 0, 5846 => 0, 5847 => 0, 5848 => 0, 5849 => 0, 5850 => 0, 5851 => 0, 5852 => 1, 5853 => 1, 5854 => 1, 5855 => 1, 5856 => 1, 5857 => 1, 5858 => 1, 5859 => 1, 5860 => 1, 5861 => 1, 5862 => 1, 5863 => 1, 5864 => 1, 5865 => 1, 5866 => 1, 5867 => 1, 5868 => 1, 5869 => 1, 5870 => 1, 5871 => 1, 5872 => 1, 5873 => 1, 5874 => 1, 5875 => 1, 5876 => 1, 5877 => 1, 5878 => 1, 5879 => 1, 5880 => 1, 5881 => 1, 5882 => 1, 5883 => 1, 5884 => 1, 5885 => 1, 5886 => 1, 5887 => 1, 5888 => 1, 5889 => 1, 5890 => 1, 5891 => 1, 5892 => 1, 5893 => 1, 5894 => 1, 5895 => 1, 5896 => 0, 5897 => 0, 5898 => 0, 5899 => 0, 5900 => 0, 5901 => 0, 5902 => 0, 5903 => 0, 5904 => 1, 5905 => 1, 5906 => 1, 5907 => 1, 5908 => 1, 5909 => 1, 5910 => 1, 5911 => 1, 5912 => 1, 5913 => 1, 5914 => 1, 5915 => 1, 5916 => 0, 5917 => 0, 5918 => 0, 5919 => 0, 5920 => 0, 5921 => 0, 5922 => 0, 5923 => 0, 5924 => 0, 5925 => 0, 5926 => 0, 5927 => 0, 5928 => 0, 5929 => 0, 5930 => 0, 5931 => 0, 5932 => 0, 5933 => 0, 5934 => 0, 
5935 => 0, 5936 => 1, 5937 => 1, 5938 => 1, 5939 => 1, 5940 => 1, 5941 => 1, 5942 => 1, 5943 => 1, 5944 => 1, 5945 => 1, 5946 => 1, 5947 => 0, 5948 => 
0, 5949 => 0, 5950 => 0, 5951 => 0, 5952 => 0, 5953 => 0, 5954 => 0, 5955 => 1, 5956 => 1, 5957 => 1, 5958 => 1, 5959 => 1, 5960 => 1, 5961 => 1, 5962 
=> 1, 5963 => 1, 5964 => 1, 5965 => 1, 5966 => 1, 5967 => 0, 5968 => 0, 5969 => 0, 5970 => 0, 5971 => 0, 5972 => 0, 5973 => 0, 5974 => 0, 5975 => 0, 5976 => 0, 5977 => 0, 5978 => 0, 5979 => 0, 5980 => 0, 5981 => 0, 5982 => 0, 5983 => 0, 5984 => 0, 5985 => 0, 5986 => 0, 5987 => 0, 5988 => 0, 5989 => 0, 5990 => 0, 5991 => 0, 5992 => 0, 5993 => 0, 5994 => 0, 5995 => 0, 5996 => 0, 5997 => 0, 5998 => 0, 5999 => 0, 6000 => 0, 6001 => 1, 6002 => 1, 6003 => 1, 6004 => 1, 6005 => 1, 6006 => 1, 6007 => 1, 6008 => 1, 6009 => 1, 6010 => 1, 6011 => 1, 6012 => 0, 6013 => 0, 6014 => 0, 6015 => 0, 6016 => 0, 6017 => 0, 6018 => 0, 6019 => 0, 6020 => 0, 6021 => 0, 6022 => 0, 6023 => 0, 6024 => 0, 6025 => 0, 6026 => 0, 6027 => 0, 6028 => 0, 6029 => 0, 6030 => 0, 6031 => 0, 6032 => 0, 6033 => 1, 6034 => 1, 6035 => 1, 6036 => 1, 6037 => 1, 6038 => 1, 6039 => 1, 6040 => 1, 6041 => 1, 6042 => 1, 6043 => 1, 6044 => 0, 6045 => 0, 6046 => 0, 6047 => 0, 6048 => 0, 6049 => 0, 6050 => 0, 6051 => 0, 6052 => 1, 6053 => 1, 6054 => 1, 6055 => 1, 6056 => 1, 6057 => 1, 6058 => 1, 6059 => 1, 6060 => 1, 6061 => 1, 6062 => 1, 6063 => 1, 6064 => 1, 6065 => 1, 6066 => 1, 6067 => 1, 6068 => 1, 6069 => 1, 6070 => 1, 6071 => 1, 6072 => 1, 6073 => 1, 6074 => 1, 6075 => 1, 6076 => 1, 6077 => 1, 6078 => 1, 6079 => 1, 6080 => 1, 6081 => 1, 6082 => 1, 6083 => 1, 6084 => 1, 6085 => 1, 
6086 => 1, 6087 => 1, 6088 => 1, 6089 => 1, 6090 => 1, 6091 => 1, 6092 => 1, 6093 => 1, 6094 => 1, 6095 => 1, 6096 => 0, 6097 => 0, 6098 => 0, 6099 => 
0, 6100 => 0, 6101 => 0, 6102 => 0, 6103 => 0, 6104 => 1, 6105 => 1, 6106 => 1, 6107 => 1, 6108 => 1, 6109 => 1, 6110 => 1, 6111 => 1, 6112 => 1, 6113 
=> 1, 6114 => 1, 6115 => 1, 6116 => 0, 6117 => 0, 6118 => 0, 6119 => 0, 6120 => 0, 6121 => 0, 6122 => 0, 6123 => 0, 6124 => 0, 6125 => 0, 6126 => 0, 6127 => 0, 6128 => 0, 6129 => 0, 6130 => 0, 6131 => 0, 6132 => 0, 6133 => 0, 6134 => 0, 6135 => 0, 6136 => 1, 6137 => 1, 6138 => 1, 6139 => 1, 6140 => 1, 6141 => 1, 6142 => 1, 6143 => 1, 6144 => 1, 6145 => 1, 6146 => 1, 6147 => 0, 6148 => 0, 6149 => 0, 6150 => 0, 6151 => 0, 6152 => 0, 6153 => 0, 6154 => 0, 6155 => 1, 6156 => 1, 6157 => 1, 6158 => 1, 6159 => 1, 6160 => 1, 6161 => 1, 6162 => 1, 6163 => 1, 6164 => 1, 6165 => 1, 6166 => 1, 6167 => 0, 6168 => 0, 6169 => 0, 6170 => 0, 6171 => 0, 6172 => 0, 6173 => 0, 6174 => 0, 6175 => 0, 6176 => 0, 6177 => 0, 6178 => 0, 6179 => 0, 6180 => 0, 6181 => 0, 6182 => 0, 6183 => 0, 6184 => 0, 6185 => 0, 6186 => 0, 6187 => 0, 6188 => 0, 6189 => 0, 6190 => 0, 6191 => 0, 6192 => 0, 6193 => 0, 6194 => 0, 6195 => 0, 6196 => 0, 6197 => 0, 6198 => 0, 6199 => 0, 6200 => 0, 6201 => 1, 6202 => 1, 6203 => 1, 6204 => 1, 6205 => 1, 6206 => 1, 6207 => 1, 6208 => 1, 6209 => 1, 6210 => 1, 6211 => 1, 6212 => 0, 6213 => 0, 6214 => 0, 6215 => 0, 6216 => 0, 6217 => 0, 6218 => 0, 6219 => 0, 6220 => 0, 6221 => 0, 6222 => 0, 6223 => 0, 6224 => 0, 6225 => 0, 6226 => 0, 6227 => 0, 6228 => 0, 6229 => 0, 6230 => 0, 6231 => 0, 6232 => 0, 6233 => 1, 6234 => 1, 6235 => 1, 6236 => 1, 
6237 => 1, 6238 => 1, 6239 => 1, 6240 => 1, 6241 => 1, 6242 => 1, 6243 => 1, 6244 => 0, 6245 => 0, 6246 => 0, 6247 => 0, 6248 => 0, 6249 => 0, 6250 => 
0, 6251 => 0, 6252 => 1, 6253 => 1, 6254 => 1, 6255 => 1, 6256 => 1, 6257 => 1, 6258 => 1, 6259 => 1, 6260 => 1, 6261 => 1, 6262 => 1, 6263 => 1, 6264 
=> 1, 6265 => 1, 6266 => 1, 6267 => 1, 6268 => 1, 6269 => 1, 6270 => 1, 6271 => 1, 6272 => 1, 6273 => 1, 6274 => 1, 6275 => 1, 6276 => 1, 6277 => 1, 6278 => 1, 6279 => 1, 6280 => 1, 6281 => 1, 6282 => 1, 6283 => 1, 6284 => 1, 6285 => 1, 6286 => 1, 6287 => 1, 6288 => 1, 6289 => 1, 6290 => 1, 6291 => 1, 6292 => 1, 6293 => 1, 6294 => 1, 6295 => 1, 6296 => 0, 6297 => 0, 6298 => 0, 6299 => 0, 6300 => 0, 6301 => 0, 6302 => 0, 6303 => 0, 6304 => 1, 6305 => 1, 6306 => 1, 6307 => 1, 6308 => 1, 6309 => 1, 6310 => 1, 6311 => 1, 6312 => 1, 6313 => 1, 6314 => 1, 6315 => 1, 6316 => 0, 6317 => 0, 6318 => 0, 6319 => 0, 6320 => 0, 6321 => 0, 6322 => 0, 6323 => 0, 6324 => 0, 6325 => 0, 6326 => 0, 6327 => 0, 6328 => 0, 6329 => 0, 6330 => 0, 6331 => 0, 6332 => 0, 6333 => 0, 6334 => 0, 6335 => 0, 6336 => 1, 6337 => 1, 6338 => 1, 6339 => 1, 6340 => 1, 6341 => 1, 6342 => 1, 6343 => 1, 6344 => 1, 6345 => 1, 6346 => 1, 6347 => 0, 6348 => 0, 6349 => 0, 6350 => 0, 6351 => 0, 6352 => 0, 6353 => 0, 6354 => 0, 6355 => 1, 6356 => 1, 6357 => 1, 6358 => 1, 6359 => 1, 6360 => 1, 6361 => 1, 6362 => 1, 6363 => 1, 6364 => 1, 6365 => 1, 6366 => 1, 6367 => 0, 6368 => 0, 6369 => 0, 6370 => 0, 6371 => 0, 6372 => 0, 6373 => 0, 6374 => 0, 6375 => 0, 6376 => 0, 6377 => 0, 6378 => 0, 6379 => 0, 6380 => 0, 6381 => 0, 6382 => 0, 6383 => 0, 6384 => 0, 6385 => 0, 6386 => 0, 6387 => 0, 
6388 => 0, 6389 => 0, 6390 => 0, 6391 => 0, 6392 => 0, 6393 => 0, 6394 => 0, 6395 => 0, 6396 => 0, 6397 => 0, 6398 => 0, 6399 => 0, 6400 => 0, 6401 => 
1, 6402 => 1, 6403 => 1, 6404 => 1, 6405 => 1, 6406 => 1, 6407 => 1, 6408 => 1, 6409 => 1, 6410 => 1, 6411 => 1, 6412 => 0, 6413 => 0, 6414 => 0, 6415 
=> 0, 6416 => 0, 6417 => 0, 6418 => 0, 6419 => 0, 6420 => 0, 6421 => 0, 6422 => 0, 6423 => 0, 6424 => 0, 6425 => 0, 6426 => 0, 6427 => 0, 6428 => 0, 6429 => 0, 6430 => 0, 6431 => 0, 6432 => 0, 6433 => 1, 6434 => 1, 6435 => 1, 6436 => 1, 6437 => 1, 6438 => 1, 6439 => 1, 6440 => 1, 6441 => 1, 6442 => 1, 6443 => 1, 6444 => 0, 6445 => 0, 6446 => 0, 6447 => 0, 6448 => 0, 6449 => 0, 6450 => 0, 6451 => 0, 6452 => 1, 6453 => 1, 6454 => 1, 6455 => 1, 6456 => 1, 6457 => 1, 6458 => 1, 6459 => 1, 6460 => 1, 6461 => 1, 6462 => 1, 6463 => 1, 6464 => 0, 6465 => 0, 6466 => 0, 6467 => 0, 6468 => 0, 6469 => 0, 6470 => 0, 6471 => 0, 6472 => 0, 6473 => 0, 6474 => 0, 6475 => 0, 6476 => 0, 6477 => 0, 6478 => 0, 6479 => 0, 6480 => 0, 6481 => 0, 6482 => 0, 6483 => 0, 6484 => 1, 6485 => 1, 6486 => 1, 6487 => 1, 6488 => 1, 6489 => 1, 6490 => 1, 6491 => 1, 6492 => 1, 6493 => 1, 6494 => 1, 6495 => 1, 6496 => 0, 6497 => 0, 6498 => 0, 6499 => 0, 6500 => 0, 6501 => 0, 6502 => 0, 6503 => 0, 6504 => 1, 6505 => 1, 6506 => 1, 6507 => 1, 6508 => 1, 6509 => 1, 6510 => 1, 6511 => 1, 6512 => 1, 6513 => 1, 6514 => 1, 6515 => 1, 6516 => 0, 6517 => 0, 6518 => 0, 6519 => 0, 6520 => 0, 6521 => 0, 6522 => 0, 6523 => 0, 6524 => 0, 6525 => 0, 6526 => 0, 6527 => 0, 6528 => 0, 6529 => 0, 6530 => 0, 6531 => 0, 6532 => 0, 6533 => 0, 6534 => 0, 6535 => 0, 6536 => 1, 6537 => 1, 6538 => 1, 
6539 => 1, 6540 => 1, 6541 => 1, 6542 => 1, 6543 => 1, 6544 => 1, 6545 => 1, 6546 => 1, 6547 => 0, 6548 => 0, 6549 => 0, 6550 => 0, 6551 => 0, 6552 => 
0, 6553 => 0, 6554 => 0, 6555 => 1, 6556 => 1, 6557 => 1, 6558 => 1, 6559 => 1, 6560 => 1, 6561 => 1, 6562 => 1, 6563 => 1, 6564 => 1, 6565 => 1, 6566 
=> 1, 6567 => 0, 6568 => 0, 6569 => 0, 6570 => 0, 6571 => 0, 6572 => 0, 6573 => 0, 6574 => 0, 6575 => 0, 6576 => 0, 6577 => 0, 6578 => 0, 6579 => 0, 6580 => 0, 6581 => 0, 6582 => 0, 6583 => 0, 6584 => 0, 6585 => 0, 6586 => 0, 6587 => 0, 6588 => 0, 6589 => 0, 6590 => 0, 6591 => 0, 6592 => 0, 6593 => 0, 6594 => 0, 6595 => 0, 6596 => 0, 6597 => 0, 6598 => 0, 6599 => 0, 6600 => 0, 6601 => 1, 6602 => 1, 6603 => 1, 6604 => 1, 6605 => 1, 6606 => 1, 6607 => 1, 6608 => 1, 6609 => 1, 6610 => 1, 6611 => 1, 6612 => 0, 6613 => 0, 6614 => 0, 6615 => 0, 6616 => 0, 6617 => 0, 6618 => 0, 6619 => 0, 6620 => 0, 6621 => 0, 6622 => 0, 6623 => 0, 6624 => 0, 6625 => 0, 6626 => 0, 6627 => 0, 6628 => 0, 6629 => 0, 6630 => 0, 6631 => 0, 6632 => 0, 6633 => 1, 6634 => 1, 6635 => 1, 6636 => 1, 6637 => 1, 6638 => 1, 6639 => 1, 6640 => 1, 6641 => 1, 6642 => 1, 6643 => 1, 6644 => 0, 6645 => 0, 6646 => 0, 6647 => 0, 6648 => 0, 6649 => 0, 6650 => 0, 6651 => 0, 6652 => 1, 6653 => 1, 6654 => 1, 6655 => 1, 6656 => 1, 6657 => 1, 6658 => 1, 6659 => 1, 6660 => 1, 6661 => 1, 6662 => 1, 6663 => 1, 6664 => 0, 6665 => 0, 6666 => 0, 6667 => 0, 6668 => 0, 6669 => 0, 6670 => 0, 6671 => 0, 6672 => 0, 6673 => 0, 6674 => 0, 6675 => 0, 6676 => 0, 6677 => 0, 6678 => 0, 6679 => 0, 6680 => 0, 6681 => 0, 6682 => 0, 6683 => 0, 6684 => 1, 6685 => 1, 6686 => 1, 6687 => 1, 6688 => 1, 6689 => 1, 
6690 => 1, 6691 => 1, 6692 => 1, 6693 => 1, 6694 => 1, 6695 => 1, 6696 => 0, 6697 => 0, 6698 => 0, 6699 => 0, 6700 => 0, 6701 => 0, 6702 => 0, 6703 => 
0, 6704 => 1, 6705 => 1, 6706 => 1, 6707 => 1, 6708 => 1, 6709 => 1, 6710 => 1, 6711 => 1, 6712 => 1, 6713 => 1, 6714 => 1, 6715 => 1, 6716 => 0, 6717 
=> 0, 6718 => 0, 6719 => 0, 6720 => 0, 6721 => 0, 6722 => 0, 6723 => 0, 6724 => 0, 6725 => 0, 6726 => 0, 6727 => 0, 6728 => 0, 6729 => 0, 6730 => 0, 6731 => 0, 6732 => 0, 6733 => 0, 6734 => 0, 6735 => 0, 6736 => 1, 6737 => 1, 6738 => 1, 6739 => 1, 6740 => 1, 6741 => 1, 6742 => 1, 6743 => 1, 6744 => 1, 6745 => 1, 6746 => 1, 6747 => 0, 6748 => 0, 6749 => 0, 6750 => 0, 6751 => 0, 6752 => 0, 6753 => 0, 6754 => 0, 6755 => 1, 6756 => 1, 6757 => 1, 6758 => 1, 6759 => 1, 6760 => 1, 6761 => 1, 6762 => 1, 6763 => 1, 6764 => 1, 6765 => 1, 6766 => 1, 6767 => 0, 6768 => 0, 6769 => 0, 6770 => 0, 6771 => 0, 6772 => 0, 6773 => 0, 6774 => 0, 6775 => 0, 6776 => 0, 6777 => 0, 6778 => 0, 6779 => 0, 6780 => 0, 6781 => 0, 6782 => 0, 6783 => 0, 6784 => 0, 6785 => 0, 6786 => 0, 6787 => 0, 6788 => 0, 6789 => 0, 6790 => 0, 6791 => 0, 6792 => 0, 6793 => 0, 6794 => 0, 6795 => 0, 6796 => 0, 6797 => 0, 6798 => 0, 6799 => 0, 6800 => 0, 6801 => 1, 6802 => 1, 6803 => 1, 6804 => 1, 6805 => 1, 6806 => 1, 6807 => 1, 6808 => 1, 6809 => 1, 6810 => 1, 6811 => 1, 6812 => 0, 6813 => 0, 6814 => 0, 6815 => 0, 6816 => 0, 6817 => 0, 6818 => 0, 6819 => 0, 6820 => 0, 6821 => 0, 6822 => 0, 6823 => 0, 6824 => 0, 6825 => 0, 6826 => 0, 6827 => 0, 6828 => 0, 6829 => 0, 6830 => 0, 6831 => 0, 6832 => 0, 6833 => 1, 6834 => 1, 6835 => 1, 6836 => 1, 6837 => 1, 6838 => 1, 6839 => 1, 6840 => 1, 
6841 => 1, 6842 => 1, 6843 => 1, 6844 => 0, 6845 => 0, 6846 => 0, 6847 => 0, 6848 => 0, 6849 => 0, 6850 => 0, 6851 => 0, 6852 => 1, 6853 => 1, 6854 => 
1, 6855 => 1, 6856 => 1, 6857 => 1, 6858 => 1, 6859 => 1, 6860 => 1, 6861 => 1, 6862 => 1, 6863 => 1, 6864 => 0, 6865 => 0, 6866 => 0, 6867 => 0, 6868 
=> 0, 6869 => 0, 6870 => 0, 6871 => 0, 6872 => 0, 6873 => 0, 6874 => 0, 6875 => 0, 6876 => 0, 6877 => 0, 6878 => 0, 6879 => 0, 6880 => 0, 6881 => 0, 6882 => 0, 6883 => 0, 6884 => 1, 6885 => 1, 6886 => 1, 6887 => 1, 6888 => 1, 6889 => 1, 6890 => 1, 6891 => 1, 6892 => 1, 6893 => 1, 6894 => 1, 6895 => 1, 6896 => 0, 6897 => 0, 6898 => 0, 6899 => 0, 6900 => 0, 6901 => 0, 6902 => 0, 6903 => 0, 6904 => 1, 6905 => 1, 6906 => 1, 6907 => 1, 6908 => 1, 6909 => 1, 6910 => 1, 6911 => 1, 6912 => 1, 6913 => 1, 6914 => 1, 6915 => 1, 6916 => 0, 6917 => 0, 6918 => 0, 6919 => 0, 6920 => 0, 6921 => 0, 6922 => 0, 6923 => 0, 6924 => 0, 6925 => 0, 6926 => 0, 6927 => 0, 6928 => 0, 6929 => 0, 6930 => 0, 6931 => 0, 6932 => 0, 6933 => 0, 6934 => 0, 6935 => 0, 6936 => 1, 6937 => 1, 6938 => 1, 6939 => 1, 6940 => 1, 6941 => 1, 6942 => 1, 6943 => 1, 6944 => 1, 6945 => 1, 6946 => 1, 6947 => 0, 6948 => 0, 6949 => 0, 6950 => 0, 6951 => 0, 6952 => 0, 6953 => 0, 6954 => 0, 6955 => 1, 6956 => 1, 6957 => 1, 6958 => 1, 6959 => 1, 6960 => 1, 6961 => 1, 6962 => 1, 6963 => 1, 6964 => 1, 6965 => 1, 6966 => 1, 6967 => 0, 6968 => 0, 6969 => 0, 6970 => 0, 6971 => 0, 6972 => 0, 6973 => 0, 6974 => 0, 6975 => 0, 6976 => 0, 6977 => 0, 6978 => 0, 6979 => 0, 6980 => 0, 6981 => 0, 6982 => 0, 6983 => 0, 6984 => 0, 6985 => 0, 6986 => 0, 6987 => 0, 6988 => 0, 6989 => 0, 6990 => 0, 6991 => 0, 
6992 => 0, 6993 => 0, 6994 => 0, 6995 => 0, 6996 => 0, 6997 => 0, 6998 => 0, 6999 => 0, 7000 => 0, 7001 => 1, 7002 => 1, 7003 => 1, 7004 => 1, 7005 => 
1, 7006 => 1, 7007 => 1, 7008 => 1, 7009 => 1, 7010 => 1, 7011 => 1, 7012 => 0, 7013 => 0, 7014 => 0, 7015 => 0, 7016 => 0, 7017 => 0, 7018 => 0, 7019 
=> 0, 7020 => 0, 7021 => 0, 7022 => 0, 7023 => 0, 7024 => 0, 7025 => 0, 7026 => 0, 7027 => 0, 7028 => 0, 7029 => 0, 7030 => 0, 7031 => 0, 7032 => 0, 7033 => 1, 7034 => 1, 7035 => 1, 7036 => 1, 7037 => 1, 7038 => 1, 7039 => 1, 7040 => 1, 7041 => 1, 7042 => 1, 7043 => 1, 7044 => 0, 7045 => 0, 7046 => 0, 7047 => 0, 7048 => 0, 7049 => 0, 7050 => 0, 7051 => 0, 7052 => 1, 7053 => 1, 7054 => 1, 7055 => 1, 7056 => 1, 7057 => 1, 7058 => 1, 7059 => 1, 7060 => 1, 7061 => 1, 7062 => 1, 7063 => 1, 7064 => 0, 7065 => 0, 7066 => 0, 7067 => 0, 7068 => 0, 7069 => 0, 7070 => 0, 7071 => 0, 7072 => 0, 7073 => 0, 7074 => 0, 7075 => 0, 7076 => 0, 7077 => 0, 7078 => 0, 7079 => 0, 7080 => 0, 7081 => 0, 7082 => 0, 7083 => 0, 7084 => 1, 7085 => 1, 7086 => 1, 7087 => 1, 7088 => 1, 7089 => 1, 7090 => 1, 7091 => 1, 7092 => 1, 7093 => 1, 7094 => 1, 7095 => 1, 7096 => 0, 7097 => 0, 7098 => 0, 7099 => 0, 7100 => 0, 7101 => 0, 7102 => 0, 7103 => 0, 7104 => 1, 7105 => 1, 7106 => 1, 7107 => 1, 7108 => 1, 7109 => 1, 7110 => 1, 7111 => 1, 7112 => 1, 7113 => 1, 7114 => 1, 7115 => 1, 7116 => 0, 7117 => 0, 7118 => 0, 7119 => 0, 7120 => 0, 7121 => 0, 7122 => 0, 7123 => 0, 7124 => 0, 7125 => 0, 7126 => 0, 7127 => 0, 7128 => 0, 7129 => 0, 7130 => 0, 7131 => 0, 7132 => 0, 7133 => 0, 7134 => 0, 7135 => 0, 7136 => 1, 7137 => 1, 7138 => 1, 7139 => 1, 7140 => 1, 7141 => 1, 7142 => 1, 
7143 => 1, 7144 => 1, 7145 => 1, 7146 => 1, 7147 => 0, 7148 => 0, 7149 => 0, 7150 => 0, 7151 => 0, 7152 => 0, 7153 => 0, 7154 => 0, 7155 => 1, 7156 => 
1, 7157 => 1, 7158 => 1, 7159 => 1, 7160 => 1, 7161 => 1, 7162 => 1, 7163 => 1, 7164 => 1, 7165 => 1, 7166 => 1, 7167 => 0, 7168 => 0, 7169 => 0, 7170 
=> 0, 7171 => 0, 7172 => 0, 7173 => 0, 7174 => 0, 7175 => 0, 7176 => 0, 7177 => 0, 7178 => 0, 7179 => 0, 7180 => 0, 7181 => 0, 7182 => 0, 7183 => 0, 7184 => 0, 7185 => 0, 7186 => 0, 7187 => 0, 7188 => 0, 7189 => 0, 7190 => 0, 7191 => 0, 7192 => 0, 7193 => 0, 7194 => 0, 7195 => 0, 7196 => 0, 7197 => 0, 7198 => 0, 7199 => 0, 7200 => 0, 7201 => 1, 7202 => 1, 7203 => 1, 7204 => 1, 7205 => 1, 7206 => 1, 7207 => 1, 7208 => 1, 7209 => 1, 7210 => 1, 7211 => 1, 7212 => 0, 7213 => 0, 7214 => 0, 7215 => 0, 7216 => 0, 7217 => 0, 7218 => 0, 7219 => 0, 7220 => 0, 7221 => 0, 7222 => 0, 7223 => 0, 7224 => 0, 7225 => 0, 7226 => 0, 7227 => 0, 7228 => 0, 7229 => 0, 7230 => 0, 7231 => 0, 7232 => 0, 7233 => 1, 7234 => 1, 7235 => 1, 7236 => 1, 7237 => 1, 7238 => 1, 7239 => 1, 7240 => 1, 7241 => 1, 7242 => 1, 7243 => 1, 7244 => 0, 7245 => 0, 7246 => 0, 7247 => 0, 7248 => 0, 7249 => 0, 7250 => 0, 7251 => 0, 7252 => 1, 7253 => 1, 7254 => 1, 7255 => 1, 7256 => 1, 7257 => 1, 7258 => 1, 7259 => 1, 7260 => 1, 7261 => 1, 7262 => 1, 7263 => 1, 7264 => 0, 7265 => 0, 7266 => 0, 7267 => 0, 7268 => 0, 7269 => 0, 7270 => 0, 7271 => 0, 7272 => 0, 7273 => 0, 7274 => 0, 7275 => 0, 7276 => 0, 7277 => 0, 7278 => 0, 7279 => 0, 7280 => 0, 7281 => 0, 7282 => 0, 7283 => 0, 7284 => 1, 7285 => 1, 7286 => 1, 7287 => 1, 7288 => 1, 7289 => 1, 7290 => 1, 7291 => 1, 7292 => 1, 7293 => 1, 
7294 => 1, 7295 => 1, 7296 => 0, 7297 => 0, 7298 => 0, 7299 => 0, 7300 => 0, 7301 => 0, 7302 => 0, 7303 => 0, 7304 => 1, 7305 => 1, 7306 => 1, 7307 => 
1, 7308 => 1, 7309 => 1, 7310 => 1, 7311 => 1, 7312 => 1, 7313 => 1, 7314 => 1, 7315 => 1, 7316 => 0, 7317 => 0, 7318 => 0, 7319 => 0, 7320 => 0, 7321 
=> 0, 7322 => 0, 7323 => 0, 7324 => 0, 7325 => 0, 7326 => 0, 7327 => 0, 7328 => 0, 7329 => 0, 7330 => 0, 7331 => 0, 7332 => 0, 7333 => 0, 7334 => 0, 7335 => 0, 7336 => 1, 7337 => 1, 7338 => 1, 7339 => 1, 7340 => 1, 7341 => 1, 7342 => 1, 7343 => 1, 7344 => 1, 7345 => 1, 7346 => 1, 7347 => 0, 7348 => 0, 7349 => 0, 7350 => 0, 7351 => 0, 7352 => 0, 7353 => 0, 7354 => 0, 7355 => 1, 7356 => 1, 7357 => 1, 7358 => 1, 7359 => 1, 7360 => 1, 7361 => 1, 7362 => 1, 7363 => 1, 7364 => 1, 7365 => 1, 7366 => 1, 7367 => 0, 7368 => 0, 7369 => 0, 7370 => 0, 7371 => 0, 7372 => 0, 7373 => 0, 7374 => 0, 7375 => 0, 7376 => 0, 7377 => 0, 7378 => 0, 7379 => 0, 7380 => 0, 7381 => 0, 7382 => 0, 7383 => 0, 7384 => 0, 7385 => 0, 7386 => 0, 7387 => 0, 7388 => 0, 7389 => 0, 7390 => 0, 7391 => 0, 7392 => 0, 7393 => 0, 7394 => 0, 7395 => 0, 7396 => 0, 7397 => 0, 7398 => 0, 7399 => 0, 7400 => 0, 7401 => 1, 7402 => 1, 7403 => 1, 7404 => 1, 7405 => 1, 7406 => 1, 7407 => 1, 7408 => 1, 7409 => 1, 7410 => 1, 7411 => 1, 7412 => 0, 7413 => 0, 7414 => 0, 7415 => 0, 7416 => 0, 7417 => 0, 7418 => 0, 7419 => 0, 7420 => 0, 7421 => 0, 7422 => 0, 7423 => 0, 7424 => 0, 7425 => 0, 7426 => 0, 7427 => 0, 7428 => 0, 7429 => 0, 7430 => 0, 7431 => 0, 7432 => 0, 7433 => 1, 7434 => 1, 7435 => 1, 7436 => 1, 7437 => 1, 7438 => 1, 7439 => 1, 7440 => 1, 7441 => 1, 7442 => 1, 7443 => 1, 7444 => 0, 
7445 => 0, 7446 => 0, 7447 => 0, 7448 => 0, 7449 => 0, 7450 => 0, 7451 => 0, 7452 => 1, 7453 => 1, 7454 => 1, 7455 => 1, 7456 => 1, 7457 => 1, 7458 => 
1, 7459 => 1, 7460 => 1, 7461 => 1, 7462 => 1, 7463 => 1, 7464 => 0, 7465 => 0, 7466 => 0, 7467 => 0, 7468 => 0, 7469 => 0, 7470 => 0, 7471 => 0, 7472 
=> 0, 7473 => 0, 7474 => 0, 7475 => 0, 7476 => 0, 7477 => 0, 7478 => 0, 7479 => 0, 7480 => 0, 7481 => 0, 7482 => 0, 7483 => 0, 7484 => 1, 7485 => 1, 7486 => 1, 7487 => 1, 7488 => 1, 7489 => 1, 7490 => 1, 7491 => 1, 7492 => 1, 7493 => 1, 7494 => 1, 7495 => 1, 7496 => 0, 7497 => 0, 7498 => 0, 7499 => 0, 7500 => 0, 7501 => 0, 7502 => 0, 7503 => 0, 7504 => 1, 7505 => 1, 7506 => 1, 7507 => 1, 7508 => 1, 7509 => 1, 7510 => 1, 7511 => 1, 7512 => 1, 7513 => 1, 7514 => 1, 7515 => 1, 7516 => 0, 7517 => 0, 7518 => 0, 7519 => 0, 7520 => 0, 7521 => 0, 7522 => 0, 7523 => 0, 7524 => 0, 7525 => 0, 7526 => 0, 7527 => 0, 7528 => 0, 7529 => 0, 7530 => 0, 7531 => 0, 7532 => 0, 7533 => 0, 7534 => 0, 7535 => 0, 7536 => 1, 7537 => 1, 7538 => 1, 7539 => 1, 7540 => 1, 7541 => 1, 7542 => 1, 7543 => 1, 7544 => 1, 7545 => 1, 7546 => 1, 7547 => 0, 7548 => 0, 7549 => 0, 7550 => 0, 7551 => 0, 7552 => 0, 7553 => 0, 7554 => 0, 7555 => 1, 7556 => 1, 7557 => 1, 7558 => 1, 7559 => 1, 7560 => 1, 7561 => 1, 7562 => 1, 7563 => 1, 7564 => 1, 7565 => 1, 7566 => 1, 7567 => 0, 7568 => 0, 7569 => 0, 7570 => 0, 7571 => 0, 7572 => 0, 7573 => 0, 7574 => 0, 7575 => 0, 7576 => 0, 7577 => 0, 7578 => 0, 7579 => 0, 7580 => 0, 7581 => 0, 7582 => 0, 7583 => 0, 7584 => 0, 7585 => 0, 7586 => 0, 7587 => 0, 7588 => 0, 7589 => 0, 7590 => 0, 7591 => 0, 7592 => 0, 7593 => 0, 7594 => 0, 7595 => 0, 
7596 => 0, 7597 => 0, 7598 => 0, 7599 => 0, 7600 => 0, 7601 => 0, 7602 => 0, 7603 => 0, 7604 => 0, 7605 => 0, 7606 => 0, 7607 => 1, 7608 => 1, 7609 => 
1, 7610 => 1, 7611 => 1, 7612 => 0, 7613 => 0, 7614 => 0, 7615 => 0, 7616 => 0, 7617 => 0, 7618 => 0, 7619 => 0, 7620 => 0, 7621 => 0, 7622 => 0, 7623 
=> 0, 7624 => 0, 7625 => 0, 7626 => 0, 7627 => 0, 7628 => 0, 7629 => 0, 7630 => 0, 7631 => 0, 7632 => 0, 7633 => 1, 7634 => 1, 7635 => 1, 7636 => 1, 7637 => 1, 7638 => 0, 7639 => 0, 7640 => 0, 7641 => 0, 7642 => 0, 7643 => 0, 7644 => 0, 7645 => 0, 7646 => 0, 7647 => 0, 7648 => 0, 7649 => 0, 7650 => 0, 7651 => 0, 7652 => 1, 7653 => 1, 7654 => 1, 7655 => 1, 7656 => 1, 7657 => 1, 7658 => 1, 7659 => 1, 7660 => 1, 7661 => 1, 7662 => 1, 7663 => 1, 7664 => 0, 7665 => 0, 7666 => 0, 7667 => 0, 7668 => 0, 7669 => 0, 7670 => 0, 7671 => 0, 7672 => 0, 7673 => 0, 7674 => 0, 7675 => 0, 7676 => 0, 7677 => 0, 7678 => 0, 7679 => 0, 7680 => 0, 7681 => 0, 7682 => 0, 7683 => 0, 7684 => 1, 7685 => 1, 7686 => 1, 7687 => 1, 7688 => 1, 7689 => 1, 7690 => 1, 7691 => 1, 7692 => 1, 7693 => 1, 7694 => 1, 7695 => 1, 7696 => 0, 7697 => 0, 7698 => 0, 7699 => 0, 7700 => 0, 7701 => 0, 7702 => 0, 7703 => 0, 7704 => 1, 7705 => 1, 7706 => 1, 7707 => 1, 7708 => 1, 7709 => 1, 7710 => 1, 7711 => 1, 7712 => 1, 7713 => 1, 7714 => 1, 7715 => 1, 7716 => 0, 7717 => 0, 7718 => 0, 7719 => 0, 7720 => 0, 7721 => 0, 7722 => 0, 7723 => 0, 7724 => 0, 7725 => 0, 7726 => 0, 7727 => 0, 7728 => 0, 7729 => 0, 7730 => 0, 7731 => 0, 7732 => 0, 7733 => 0, 7734 => 0, 7735 => 0, 7736 => 1, 7737 => 1, 7738 => 1, 7739 => 1, 7740 => 1, 7741 => 1, 7742 => 1, 7743 => 1, 7744 => 1, 7745 => 1, 7746 => 1, 
7747 => 0, 7748 => 0, 7749 => 0, 7750 => 0, 7751 => 0, 7752 => 0, 7753 => 0, 7754 => 0, 7755 => 1, 7756 => 1, 7757 => 1, 7758 => 1, 7759 => 1, 7760 => 
1, 7761 => 1, 7762 => 1, 7763 => 1, 7764 => 1, 7765 => 1, 7766 => 1, 7767 => 0, 7768 => 0, 7769 => 0, 7770 => 0, 7771 => 0, 7772 => 0, 7773 => 0, 7774 
=> 0, 7775 => 0, 7776 => 0, 7777 => 0, 7778 => 0, 7779 => 0, 7780 => 0, 7781 => 0, 7782 => 0, 7783 => 0, 7784 => 0, 7785 => 0, 7786 => 0, 7787 => 0, 7788 => 0, 7789 => 0, 7790 => 0, 7791 => 0, 7792 => 0, 7793 => 0, 7794 => 0, 7795 => 0, 7796 => 0, 7797 => 0, 7798 => 0, 7799 => 0, 7800 => 0, 7801 => 0, 7802 => 0, 7803 => 0, 7804 => 0, 7805 => 0, 7806 => 0, 7807 => 1, 7808 => 1, 7809 => 1, 7810 => 1, 7811 => 1, 7812 => 1, 7813 => 1, 7814 => 1, 7815 => 1, 7816 => 1, 7817 => 1, 7818 => 1, 7819 => 1, 7820 => 1, 7821 => 1, 7822 => 1, 7823 => 1, 7824 => 1, 7825 => 1, 7826 => 1, 7827 => 1, 7828 => 1, 7829 => 1, 7830 => 1, 7831 => 1, 7832 => 1, 7833 => 1, 7834 => 1, 7835 => 1, 7836 => 1, 7837 => 1, 7838 => 0, 7839 => 0, 7840 => 0, 7841 => 0, 7842 => 0, 7843 => 0, 7844 => 0, 7845 => 0, 7846 => 0, 7847 => 0, 7848 => 0, 7849 => 0, 7850 => 0, 7851 => 0, 7852 => 1, 7853 => 1, 7854 => 1, 7855 => 1, 7856 => 1, 7857 => 1, 7858 => 1, 7859 => 1, 7860 => 1, 7861 => 1, 7862 => 1, 7863 => 1, 7864 => 0, 7865 => 0, 7866 => 0, 7867 => 0, 7868 => 0, 7869 => 0, 7870 => 0, 7871 => 0, 7872 => 0, 7873 => 0, 7874 => 0, 7875 => 0, 7876 => 0, 7877 => 0, 7878 => 0, 7879 => 0, 7880 => 0, 7881 => 0, 7882 => 0, 7883 => 0, 7884 => 1, 7885 => 1, 7886 => 1, 7887 => 1, 7888 => 1, 7889 => 1, 7890 => 1, 7891 => 1, 7892 => 1, 7893 => 1, 7894 => 1, 7895 => 1, 7896 => 0, 7897 => 0, 
7898 => 0, 7899 => 0, 7900 => 0, 7901 => 0, 7902 => 0, 7903 => 0, 7904 => 1, 7905 => 1, 7906 => 1, 7907 => 1, 7908 => 1, 7909 => 1, 7910 => 1, 7911 => 
1, 7912 => 1, 7913 => 1, 7914 => 1, 7915 => 1, 7916 => 0, 7917 => 0, 7918 => 0, 7919 => 0, 7920 => 0, 7921 => 0, 7922 => 0, 7923 => 0, 7924 => 0, 7925 
=> 0, 7926 => 0, 7927 => 0, 7928 => 0, 7929 => 0, 7930 => 0, 7931 => 0, 7932 => 0, 7933 => 0, 7934 => 0, 7935 => 0, 7936 => 1, 7937 => 1, 7938 => 1, 7939 => 1, 7940 => 1, 7941 => 1, 7942 => 1, 7943 => 1, 7944 => 1, 7945 => 1, 7946 => 1, 7947 => 0, 7948 => 0, 7949 => 0, 7950 => 0, 7951 => 0, 7952 => 0, 7953 => 0, 7954 => 0, 7955 => 1, 7956 => 1, 7957 => 1, 7958 => 1, 7959 => 1, 7960 => 1, 7961 => 1, 7962 => 1, 7963 => 1, 7964 => 1, 7965 => 1, 7966 => 1, 7967 => 1, 7968 => 1, 7969 => 1, 7970 => 1, 7971 => 1, 7972 => 1, 7973 => 1, 7974 => 1, 7975 => 1, 7976 => 1, 7977 => 1, 7978 => 1, 7979 => 1, 7980 => 1, 7981 => 1, 7982 => 1, 7983 => 1, 7984 => 1, 7985 => 1, 7986 => 1, 7987 => 1, 7988 => 1, 7989 => 1, 7990 => 1, 7991 => 1, 7992 => 1, 7993 => 1, 7994 => 1, 7995 => 1, 7996 => 1, 7997 => 1, 7998 => 1, 7999 => 0, 8000 => 0, 8001 => 0, 8002 => 0, 8003 => 0, 8004 => 0, 8005 => 0, 8006 => 0, 8007 => 1, 8008 => 1, 8009 => 1, 8010 => 1, 8011 => 1, 8012 => 1, 8013 => 1, 8014 => 1, 8015 => 1, 8016 => 1, 8017 => 1, 8018 => 1, 8019 => 1, 8020 => 1, 8021 => 1, 8022 => 1, 8023 => 1, 8024 => 1, 8025 => 1, 8026 => 1, 8027 => 1, 8028 => 1, 8029 => 1, 8030 => 1, 8031 => 1, 8032 => 1, 8033 => 1, 8034 => 1, 8035 => 1, 8036 => 1, 8037 => 1, 8038 => 0, 8039 => 0, 8040 => 0, 8041 => 0, 8042 => 0, 8043 => 0, 8044 => 0, 8045 => 0, 8046 => 0, 8047 => 0, 8048 => 0, 
8049 => 0, 8050 => 0, 8051 => 0, 8052 => 1, 8053 => 1, 8054 => 1, 8055 => 1, 8056 => 1, 8057 => 1, 8058 => 1, 8059 => 1, 8060 => 1, 8061 => 1, 8062 => 
1, 8063 => 1, 8064 => 0, 8065 => 0, 8066 => 0, 8067 => 0, 8068 => 0, 8069 => 0, 8070 => 0, 8071 => 0, 8072 => 0, 8073 => 0, 8074 => 0, 8075 => 0, 8076 
=> 0, 8077 => 0, 8078 => 0, 8079 => 0, 8080 => 0, 8081 => 0, 8082 => 0, 8083 => 0, 8084 => 1, 8085 => 1, 8086 => 1, 8087 => 1, 8088 => 1, 8089 => 1, 8090 => 1, 8091 => 1, 8092 => 1, 8093 => 1, 8094 => 1, 8095 => 1, 8096 => 0, 8097 => 0, 8098 => 0, 8099 => 0, 8100 => 0, 8101 => 0, 8102 => 0, 8103 => 0, 8104 => 1, 8105 => 1, 8106 => 1, 8107 => 1, 8108 => 1, 8109 => 1, 8110 => 1, 8111 => 1, 8112 => 1, 8113 => 1, 8114 => 1, 8115 => 1, 8116 => 0, 8117 => 0, 8118 => 0, 8119 => 0, 8120 => 0, 8121 => 0, 8122 => 0, 8123 => 0, 8124 => 0, 8125 => 0, 8126 => 0, 8127 => 0, 8128 => 0, 8129 => 0, 8130 => 0, 8131 => 0, 8132 => 0, 8133 => 0, 8134 => 0, 8135 => 0, 8136 => 1, 8137 => 1, 8138 => 1, 8139 => 1, 8140 => 1, 8141 => 1, 8142 => 1, 8143 => 1, 8144 => 1, 8145 => 1, 8146 => 1, 8147 => 0, 8148 => 0, 8149 => 0, 8150 => 0, 8151 => 0, 8152 => 0, 8153 => 0, 8154 => 0, 8155 => 1, 8156 => 1, 8157 => 1, 8158 => 1, 8159 => 1, 8160 => 1, 8161 => 1, 8162 => 1, 8163 => 1, 8164 => 1, 8165 => 1, 8166 => 1, 8167 => 1, 8168 => 1, 8169 => 1, 8170 => 1, 8171 => 1, 8172 => 1, 8173 => 1, 8174 => 1, 8175 => 1, 8176 => 1, 8177 => 1, 8178 => 1, 8179 => 1, 8180 => 1, 8181 => 1, 8182 => 1, 8183 => 1, 8184 => 1, 8185 => 1, 8186 => 1, 8187 => 1, 8188 => 1, 8189 => 1, 8190 => 1, 8191 => 1, 8192 => 1, 8193 => 1, 8194 => 1, 8195 => 1, 8196 => 1, 8197 => 1, 8198 => 1, 8199 => 0, 
8200 => 0, 8201 => 0, 8202 => 0, 8203 => 0, 8204 => 0, 8205 => 0, 8206 => 0, 8207 => 1, 8208 => 1, 8209 => 1, 8210 => 1, 8211 => 1, 8212 => 1, 8213 => 
1, 8214 => 1, 8215 => 1, 8216 => 1, 8217 => 1, 8218 => 1, 8219 => 1, 8220 => 1, 8221 => 1, 8222 => 1, 8223 => 1, 8224 => 1, 8225 => 1, 8226 => 1, 8227 
=> 1, 8228 => 1, 8229 => 1, 8230 => 1, 8231 => 1, 8232 => 1, 8233 => 1, 8234 => 1, 8235 => 1, 8236 => 1, 8237 => 1, 8238 => 0, 8239 => 0, 8240 => 0, 8241 => 0, 8242 => 0, 8243 => 0, 8244 => 0, 8245 => 0, 8246 => 0, 8247 => 0, 8248 => 0, 8249 => 0, 8250 => 0, 8251 => 0, 8252 => 1, 8253 => 1, 8254 => 1, 8255 => 1, 8256 => 1, 8257 => 1, 8258 => 1, 8259 => 1, 8260 => 1, 8261 => 1, 8262 => 1, 8263 => 1, 8264 => 0, 8265 => 0, 8266 => 0, 8267 => 0, 8268 => 0, 8269 => 0, 8270 => 0, 8271 => 0, 8272 => 0, 8273 => 0, 8274 => 0, 8275 => 0, 8276 => 0, 8277 => 0, 8278 => 0, 8279 => 0, 8280 => 0, 8281 => 0, 8282 => 0, 8283 => 0, 8284 => 1, 8285 => 1, 8286 => 1, 8287 => 1, 8288 => 1, 8289 => 1, 8290 => 1, 8291 => 1, 8292 => 1, 8293 => 1, 8294 => 1, 8295 => 1, 8296 => 0, 8297 => 0, 8298 => 0, 8299 => 0, 8300 => 0, 8301 => 0, 8302 => 0, 8303 => 0, 8304 => 1, 8305 => 1, 8306 => 1, 8307 => 1, 8308 => 1, 8309 => 1, 8310 => 1, 8311 => 1, 8312 => 1, 8313 => 1, 8314 => 1, 8315 => 1, 8316 => 0, 8317 => 0, 8318 => 0, 8319 => 0, 8320 => 0, 8321 => 0, 8322 => 0, 8323 => 0, 8324 => 0, 8325 => 0, 8326 => 0, 8327 => 0, 8328 => 0, 8329 => 0, 8330 => 0, 8331 => 0, 8332 => 0, 8333 => 0, 8334 => 0, 8335 => 0, 8336 => 1, 8337 => 1, 8338 => 1, 8339 => 1, 8340 => 1, 8341 => 1, 8342 => 1, 8343 => 1, 8344 => 1, 8345 => 1, 8346 => 1, 8347 => 0, 8348 => 0, 8349 => 0, 8350 => 0, 
8351 => 0, 8352 => 0, 8353 => 0, 8354 => 0, 8355 => 1, 8356 => 1, 8357 => 1, 8358 => 1, 8359 => 1, 8360 => 1, 8361 => 1, 8362 => 1, 8363 => 1, 8364 => 
1, 8365 => 1, 8366 => 1, 8367 => 1, 8368 => 1, 8369 => 1, 8370 => 1, 8371 => 1, 8372 => 1, 8373 => 1, 8374 => 1, 8375 => 1, 8376 => 1, 8377 => 1, 8378 
=> 1, 8379 => 1, 8380 => 1, 8381 => 1, 8382 => 1, 8383 => 1, 8384 => 1, 8385 => 1, 8386 => 1, 8387 => 1, 8388 => 1, 8389 => 1, 8390 => 1, 8391 => 1, 8392 => 1, 8393 => 1, 8394 => 1, 8395 => 1, 8396 => 1, 8397 => 1, 8398 => 1, 8399 => 0, 8400 => 0, 8401 => 0, 8402 => 0, 8403 => 0, 8404 => 0, 8405 => 0, 8406 => 0, 8407 => 1, 8408 => 1, 8409 => 1, 8410 => 1, 8411 => 1, 8412 => 1, 8413 => 1, 8414 => 1, 8415 => 1, 8416 => 1, 8417 => 1, 8418 => 1, 8419 => 1, 8420 => 1, 8421 => 1, 8422 => 1, 8423 => 1, 8424 => 1, 8425 => 1, 8426 => 1, 8427 => 1, 8428 => 1, 8429 => 1, 8430 => 1, 8431 => 1, 8432 => 1, 8433 => 1, 8434 => 1, 8435 => 1, 8436 => 1, 8437 => 1, 8438 => 0, 8439 => 0, 8440 => 0, 8441 => 0, 8442 => 0, 8443 => 0, 8444 => 0, 8445 => 0, 8446 => 0, 8447 => 0, 8448 => 0, 8449 => 0, 8450 => 0, 8451 => 0, 8452 => 1, 8453 => 1, 8454 => 1, 8455 => 1, 8456 => 1, 8457 => 1, 8458 => 1, 8459 => 1, 8460 => 1, 8461 => 1, 8462 => 1, 8463 => 1, 8464 => 0, 8465 => 0, 8466 => 0, 8467 => 0, 8468 => 0, 8469 => 0, 8470 => 0, 8471 => 0, 8472 => 0, 8473 => 0, 8474 => 0, 8475 => 0, 8476 => 0, 8477 => 0, 8478 => 0, 8479 => 0, 8480 => 0, 8481 => 0, 8482 => 0, 8483 => 0, 8484 => 1, 8485 => 1, 8486 => 1, 8487 => 1, 8488 => 1, 8489 => 1, 8490 => 1, 8491 => 1, 8492 => 1, 8493 => 1, 8494 => 1, 8495 => 1, 8496 => 0, 8497 => 0, 8498 => 0, 8499 => 0, 8500 => 0, 8501 => 0, 
8502 => 0, 8503 => 0, 8504 => 1, 8505 => 1, 8506 => 1, 8507 => 1, 8508 => 1, 8509 => 1, 8510 => 1, 8511 => 1, 8512 => 1, 8513 => 1, 8514 => 1, 8515 => 
1, 8516 => 0, 8517 => 0, 8518 => 0, 8519 => 0, 8520 => 0, 8521 => 0, 8522 => 0, 8523 => 0, 8524 => 0, 8525 => 0, 8526 => 0, 8527 => 0, 8528 => 0, 8529 
=> 0, 8530 => 0, 8531 => 0, 8532 => 0, 8533 => 0, 8534 => 0, 8535 => 0, 8536 => 1, 8537 => 1, 8538 => 1, 8539 => 1, 8540 => 1, 8541 => 1, 8542 => 1, 8543 => 1, 8544 => 1, 8545 => 1, 8546 => 1, 8547 => 0, 8548 => 0, 8549 => 0, 8550 => 0, 8551 => 0, 8552 => 0, 8553 => 0, 8554 => 0, 8555 => 1, 8556 => 1, 8557 => 1, 8558 => 1, 8559 => 1, 8560 => 1, 8561 => 1, 8562 => 1, 8563 => 1, 8564 => 1, 8565 => 1, 8566 => 1, 8567 => 1, 8568 => 1, 8569 => 1, 8570 => 1, 8571 => 1, 8572 => 1, 8573 => 1, 8574 => 1, 8575 => 1, 8576 => 1, 8577 => 1, 8578 => 1, 8579 => 1, 8580 => 1, 8581 => 1, 8582 => 1, 8583 => 1, 8584 => 1, 8585 => 1, 8586 => 1, 8587 => 1, 8588 => 1, 8589 => 1, 8590 => 1, 8591 => 1, 8592 => 1, 8593 => 1, 8594 => 1, 8595 => 1, 8596 => 1, 8597 => 1, 8598 => 1, 8599 => 0, 8600 => 0, 8601 => 0, 8602 => 0, 8603 => 0, 8604 => 0, 8605 => 0, 8606 => 0, 8607 => 1, 8608 => 1, 8609 => 1, 8610 => 1, 8611 => 1, 8612 => 1, 8613 => 1, 8614 => 1, 8615 => 1, 8616 => 1, 8617 => 1, 8618 => 1, 8619 => 1, 8620 => 1, 8621 => 1, 8622 => 1, 8623 => 1, 8624 => 1, 8625 => 1, 8626 => 1, 8627 => 1, 8628 => 1, 8629 => 1, 8630 => 1, 8631 => 1, 8632 => 1, 8633 => 1, 8634 => 1, 8635 => 1, 8636 => 1, 8637 => 1, 8638 => 0, 8639 => 0, 8640 => 0, 8641 => 0, 8642 => 0, 8643 => 0, 8644 => 0, 8645 => 0, 8646 => 0, 8647 => 0, 8648 => 0, 8649 => 0, 8650 => 0, 8651 => 0, 8652 => 1, 
8653 => 1, 8654 => 1, 8655 => 1, 8656 => 1, 8657 => 1, 8658 => 1, 8659 => 1, 8660 => 1, 8661 => 1, 8662 => 1, 8663 => 1, 8664 => 0, 8665 => 0, 8666 => 
0, 8667 => 0, 8668 => 0, 8669 => 0, 8670 => 0, 8671 => 0, 8672 => 0, 8673 => 0, 8674 => 0, 8675 => 0, 8676 => 0, 8677 => 0, 8678 => 0, 8679 => 0, 8680 
=> 0, 8681 => 0, 8682 => 0, 8683 => 0, 8684 => 1, 8685 => 1, 8686 => 1, 8687 => 1, 8688 => 1, 8689 => 1, 8690 => 1, 8691 => 1, 8692 => 1, 8693 => 1, 8694 => 1, 8695 => 1, 8696 => 0, 8697 => 0, 8698 => 0, 8699 => 0, 8700 => 0, 8701 => 0, 8702 => 0, 8703 => 0, 8704 => 1, 8705 => 1, 8706 => 1, 8707 => 1, 8708 => 1, 8709 => 1, 8710 => 1, 8711 => 1, 8712 => 1, 8713 => 1, 8714 => 1, 8715 => 1, 8716 => 0, 8717 => 0, 8718 => 0, 8719 => 0, 8720 => 0, 8721 => 0, 8722 => 0, 8723 => 0, 8724 => 0, 8725 => 0, 8726 => 0, 8727 => 0, 8728 => 0, 8729 => 0, 8730 => 0, 8731 => 0, 8732 => 0, 8733 => 0, 8734 => 0, 8735 => 0, 8736 => 1, 8737 => 1, 8738 => 1, 8739 => 1, 8740 => 1, 8741 => 1, 8742 => 1, 8743 => 1, 8744 => 1, 8745 => 1, 8746 => 1, 8747 => 0, 8748 => 0, 8749 => 0, 8750 => 0, 8751 => 0, 8752 => 0, 8753 => 0, 8754 => 0, 8755 => 1, 8756 => 1, 8757 => 1, 8758 => 1, 8759 => 1, 8760 => 1, 8761 => 1, 8762 => 1, 8763 => 1, 8764 => 1, 8765 => 1, 8766 => 1, 8767 => 1, 8768 => 1, 8769 => 1, 8770 => 1, 8771 => 1, 8772 => 1, 8773 => 1, 8774 => 1, 8775 => 1, 8776 => 1, 8777 => 1, 8778 => 1, 8779 => 1, 8780 => 1, 8781 => 1, 8782 => 1, 8783 => 1, 8784 => 1, 8785 => 1, 8786 => 1, 8787 => 1, 8788 => 1, 8789 => 1, 8790 => 1, 8791 => 1, 8792 => 1, 8793 => 1, 8794 => 1, 8795 => 1, 8796 => 1, 8797 => 1, 8798 => 1, 8799 => 0, 8800 => 0, 8801 => 0, 8802 => 0, 8803 => 0, 
8804 => 0, 8805 => 0, 8806 => 0, 8807 => 1, 8808 => 1, 8809 => 1, 8810 => 1, 8811 => 1, 8812 => 1, 8813 => 1, 8814 => 1, 8815 => 1, 8816 => 1, 8817 => 
1, 8818 => 1, 8819 => 1, 8820 => 1, 8821 => 1, 8822 => 1, 8823 => 1, 8824 => 1, 8825 => 1, 8826 => 1, 8827 => 1, 8828 => 1, 8829 => 1, 8830 => 1, 8831 
=> 1, 8832 => 1, 8833 => 1, 8834 => 1, 8835 => 1, 8836 => 1, 8837 => 1, 8838 => 0, 8839 => 0, 8840 => 0, 8841 => 0, 8842 => 0, 8843 => 0, 8844 => 0, 8845 => 0, 8846 => 0, 8847 => 0, 8848 => 0, 8849 => 0, 8850 => 0, 8851 => 0, 8852 => 1, 8853 => 1, 8854 => 1, 8855 => 1, 8856 => 1, 8857 => 1, 8858 => 1, 8859 => 1, 8860 => 1, 8861 => 1, 8862 => 1, 8863 => 1, 8864 => 0, 8865 => 0, 8866 => 0, 8867 => 0, 8868 => 0, 8869 => 0, 8870 => 0, 8871 => 0, 8872 => 0, 8873 => 0, 8874 => 0, 8875 => 0, 8876 => 0, 8877 => 0, 8878 => 0, 8879 => 0, 8880 => 0, 8881 => 0, 8882 => 0, 8883 => 0, 8884 => 1, 8885 => 1, 8886 => 1, 8887 => 1, 8888 => 1, 8889 => 1, 8890 => 1, 8891 => 1, 8892 => 1, 8893 => 1, 8894 => 1, 8895 => 1, 8896 => 0, 8897 => 0, 8898 => 0, 8899 => 0, 8900 => 0, 8901 => 0, 8902 => 0, 8903 => 0, 8904 => 1, 8905 => 1, 8906 => 1, 8907 => 1, 8908 => 1, 8909 => 1, 8910 => 1, 8911 => 1, 8912 => 1, 8913 => 1, 8914 => 1, 8915 => 1, 8916 => 0, 8917 => 0, 8918 => 0, 8919 => 0, 8920 => 0, 8921 => 0, 8922 => 0, 8923 => 0, 8924 => 0, 8925 => 0, 8926 => 0, 8927 => 0, 8928 => 0, 8929 => 0, 8930 => 0, 8931 => 0, 8932 => 0, 8933 => 0, 8934 => 0, 8935 => 0, 8936 => 1, 8937 => 1, 8938 => 1, 8939 => 1, 8940 => 1, 8941 => 1, 8942 => 1, 8943 => 1, 8944 => 1, 8945 => 1, 8946 => 1, 8947 => 0, 8948 => 0, 8949 => 0, 8950 => 0, 8951 => 0, 8952 => 0, 8953 => 0, 8954 => 0, 
8955 => 1, 8956 => 1, 8957 => 1, 8958 => 1, 8959 => 1, 8960 => 1, 8961 => 1, 8962 => 1, 8963 => 1, 8964 => 1, 8965 => 1, 8966 => 1, 8967 => 1, 8968 => 
1, 8969 => 1, 8970 => 1, 8971 => 1, 8972 => 1, 8973 => 1, 8974 => 1, 8975 => 1, 8976 => 1, 8977 => 1, 8978 => 1, 8979 => 1, 8980 => 1, 8981 => 1, 8982 
=> 1, 8983 => 1, 8984 => 1, 8985 => 1, 8986 => 1, 8987 => 1, 8988 => 1, 8989 => 1, 8990 => 1, 8991 => 1, 8992 => 1, 8993 => 1, 8994 => 1, 8995 => 1, 8996 => 1, 8997 => 1, 8998 => 1, 8999 => 0
	
	);
	
		constant rom_option_1 : rom_bitmap := (
0 => 0, 1 => 0, 2 => 0, 3 => 0, 4 => 0, 5 => 0, 6 => 0, 7 => 0, 8 => 0, 9 => 0, 10 => 0, 11 => 0, 12 => 0, 13 => 0, 14 => 0, 15 => 0, 16 => 0, 17 => 0, 18 => 0, 19 => 0, 20 => 0, 21 => 0, 22 => 0, 23 => 0, 24 => 0, 25 => 0, 26 => 0, 27 => 0, 28 => 0, 29 => 0, 30 => 0, 31 => 0, 32 => 0, 33 => 0, 34 => 
0, 35 => 0, 36 => 0, 37 => 0, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 0, 45 => 0, 46 => 0, 47 => 0, 48 => 0, 49 => 0, 50 => 0, 51 => 0, 52 => 0, 53 => 0, 54 => 0, 55 => 0, 56 => 0, 57 => 0, 58 => 0, 59 => 0, 60 => 0, 61 => 0, 62 => 0, 63 => 0, 64 => 0, 65 => 0, 66 => 0, 67 => 0, 68 => 0, 69 => 0, 70 => 0, 71 => 0, 72 => 0, 73 => 0, 74 => 0, 75 => 0, 76 => 0, 77 => 0, 78 => 0, 79 => 0, 80 => 0, 81 => 0, 82 => 0, 83 => 0, 84 => 0, 
85 => 0, 86 => 0, 87 => 0, 88 => 0, 89 => 0, 90 => 0, 91 => 0, 92 => 0, 93 => 0, 94 => 0, 95 => 0, 96 => 0, 97 => 0, 98 => 0, 99 => 0, 100 => 0, 101 => 0, 102 => 0, 103 => 0, 104 => 0, 105 => 0, 106 => 0, 107 => 0, 108 => 0, 109 => 0, 110 => 0, 111 => 0, 112 => 0, 113 => 0, 114 => 0, 115 => 0, 116 => 
0, 117 => 0, 118 => 0, 119 => 0, 120 => 0, 121 => 0, 122 => 0, 123 => 0, 124 => 0, 125 => 0, 126 => 0, 127 => 0, 128 => 0, 129 => 0, 130 => 0, 131 => 0, 132 => 0, 133 => 0, 134 => 0, 135 => 0, 136 => 0, 137 => 0, 138 => 0, 139 => 0, 140 => 0, 141 => 0, 142 => 0, 143 => 0, 144 => 0, 145 => 0, 146 => 0, 147 => 0, 148 => 0, 149 => 0, 150 => 0, 151 => 0, 152 => 0, 153 => 0, 154 => 0, 155 => 0, 156 => 0, 157 => 0, 158 => 0, 159 => 0, 160 => 0, 161 => 0, 
162 => 0, 163 => 0, 164 => 0, 165 => 0, 166 => 0, 167 => 0, 168 => 0, 169 => 0, 170 => 0, 171 => 0, 172 => 0, 173 => 0, 174 => 0, 175 => 0, 176 => 0, 177 => 0, 178 => 0, 179 => 0, 180 => 0, 181 => 0, 182 => 0, 183 => 0, 184 => 0, 185 => 0, 186 => 0, 187 => 0, 188 => 0, 189 => 0, 190 => 0, 191 => 0, 192 => 0, 193 => 0, 194 => 0, 195 => 0, 196 => 0, 197 => 0, 198 => 0, 199 => 0, 200 => 0, 201 => 0, 202 => 0, 203 => 0, 204 => 0, 205 => 0, 206 => 0, 207 => 0, 208 => 0, 209 => 0, 210 => 0, 211 => 0, 212 => 0, 213 => 0, 214 => 0, 215 => 0, 216 => 0, 217 => 0, 218 => 0, 219 => 0, 220 => 0, 221 => 0, 222 
=> 0, 223 => 0, 224 => 0, 225 => 0, 226 => 0, 227 => 0, 228 => 0, 229 => 0, 230 => 0, 231 => 0, 232 => 0, 233 => 0, 234 => 0, 235 => 0, 236 => 0, 237 => 0, 238 => 0, 239 => 0, 240 => 0, 241 => 0, 242 => 0, 243 => 0, 244 => 0, 245 => 0, 246 => 0, 247 => 1, 248 => 1, 249 => 1, 250 => 0, 251 => 0, 252 => 0, 253 => 0, 254 => 0, 255 => 0, 256 => 0, 257 => 0, 258 => 0, 259 => 0, 260 => 0, 261 => 0, 262 => 0, 263 => 0, 264 => 0, 265 => 0, 266 => 0, 267 => 
0, 268 => 0, 269 => 0, 270 => 0, 271 => 0, 272 => 0, 273 => 0, 274 => 0, 275 => 0, 276 => 0, 277 => 0, 278 => 0, 279 => 0, 280 => 0, 281 => 0, 282 => 0, 283 => 0, 284 => 0, 285 => 0, 286 => 0, 287 => 0, 288 => 0, 289 => 0, 290 => 0, 291 => 0, 292 => 0, 293 => 0, 294 => 0, 295 => 0, 296 => 0, 297 => 0, 298 => 0, 299 => 0, 300 => 0, 301 => 0, 302 => 0, 303 => 0, 304 => 0, 305 => 0, 306 => 0, 307 => 0, 308 => 0, 309 => 0, 310 => 0, 311 => 0, 312 => 0, 
313 => 0, 314 => 0, 315 => 0, 316 => 0, 317 => 0, 318 => 0, 319 => 0, 320 => 0, 321 => 0, 322 => 0, 323 => 0, 324 => 0, 325 => 0, 326 => 0, 327 => 0, 328 => 0, 329 => 0, 330 => 0, 331 => 0, 332 => 0, 333 => 0, 334 => 0, 335 => 0, 336 => 0, 337 => 0, 338 => 0, 339 => 0, 340 => 0, 341 => 0, 342 => 0, 343 => 0, 344 => 0, 345 => 0, 346 => 0, 347 => 0, 348 => 0, 349 => 0, 350 => 0, 351 => 0, 352 => 0, 353 => 0, 354 => 0, 355 => 0, 356 => 0, 357 => 0, 358 => 0, 359 => 0, 360 => 0, 361 => 0, 362 => 0, 363 => 0, 364 => 0, 365 => 0, 366 => 0, 367 => 0, 368 => 0, 369 => 0, 370 => 0, 371 => 0, 372 => 0, 373 
=> 0, 374 => 0, 375 => 0, 376 => 0, 377 => 0, 378 => 0, 379 => 0, 380 => 0, 381 => 0, 382 => 0, 383 => 0, 384 => 0, 385 => 0, 386 => 0, 387 => 0, 388 => 0, 389 => 0, 390 => 0, 391 => 0, 392 => 0, 393 => 0, 394 => 0, 395 => 0, 396 => 0, 397 => 0, 398 => 0, 399 => 0, 400 => 0, 401 => 0, 402 => 0, 403 => 0, 404 => 0, 405 => 0, 406 => 0, 407 => 0, 408 => 0, 409 => 0, 410 => 0, 411 => 1, 412 => 1, 413 => 1, 414 => 0, 415 => 0, 416 => 0, 417 => 0, 418 => 
0, 419 => 0, 420 => 0, 421 => 0, 422 => 0, 423 => 0, 424 => 0, 425 => 0, 426 => 0, 427 => 0, 428 => 0, 429 => 0, 430 => 0, 431 => 0, 432 => 0, 433 => 0, 434 => 0, 435 => 0, 436 => 0, 437 => 0, 438 => 0, 439 => 0, 440 => 0, 441 => 0, 442 => 0, 443 => 0, 444 => 0, 445 => 0, 446 => 0, 447 => 0, 448 => 0, 449 => 0, 450 => 0, 451 => 0, 452 => 0, 453 => 0, 454 => 0, 455 => 0, 456 => 0, 457 => 0, 458 => 0, 459 => 0, 460 => 0, 461 => 0, 462 => 0, 463 => 0, 
464 => 0, 465 => 0, 466 => 0, 467 => 0, 468 => 0, 469 => 0, 470 => 0, 471 => 0, 472 => 0, 473 => 0, 474 => 0, 475 => 0, 476 => 0, 477 => 0, 478 => 0, 479 => 0, 480 => 0, 481 => 0, 482 => 0, 483 => 0, 484 => 0, 485 => 0, 486 => 0, 487 => 0, 488 => 0, 489 => 0, 490 => 0, 491 => 0, 492 => 0, 493 => 0, 494 => 0, 495 => 1, 496 => 0, 497 => 0, 498 => 0, 499 => 0, 500 => 0, 501 => 0, 502 => 0, 503 => 0, 504 => 1, 505 => 0, 506 => 0, 507 => 0, 508 => 0, 509 => 0, 510 => 0, 511 => 1, 512 => 0, 513 => 0, 514 => 0, 515 => 0, 516 => 0, 517 => 0, 518 => 0, 519 => 0, 520 => 0, 521 => 0, 522 => 0, 523 => 1, 524 
=> 0, 525 => 0, 526 => 0, 527 => 0, 528 => 0, 529 => 0, 530 => 0, 531 => 0, 532 => 0, 533 => 0, 534 => 0, 535 => 0, 536 => 0, 537 => 0, 538 => 0, 539 => 0, 540 => 0, 541 => 0, 542 => 1, 543 => 0, 544 => 0, 545 => 0, 546 => 0, 547 => 0, 548 => 0, 549 => 0, 550 => 0, 551 => 0, 552 => 0, 553 => 0, 554 => 0, 555 => 0, 556 => 0, 557 => 0, 558 => 0, 559 => 0, 560 => 0, 561 => 0, 562 => 0, 563 => 0, 564 => 0, 565 => 0, 566 => 0, 567 => 0, 568 => 0, 569 => 
0, 570 => 0, 571 => 0, 572 => 0, 573 => 0, 574 => 0, 575 => 1, 576 => 1, 577 => 1, 578 => 0, 579 => 0, 580 => 0, 581 => 0, 582 => 0, 583 => 0, 584 => 1, 585 => 0, 586 => 0, 587 => 0, 588 => 0, 589 => 0, 590 => 0, 591 => 0, 592 => 0, 593 => 1, 594 => 0, 595 => 0, 596 => 0, 597 => 0, 598 => 0, 599 => 0, 600 => 0, 601 => 1, 602 => 0, 603 => 1, 604 => 0, 605 => 0, 606 => 0, 607 => 0, 608 => 0, 609 => 0, 610 => 0, 611 => 0, 612 => 0, 613 => 0, 614 => 0, 
615 => 1, 616 => 0, 617 => 0, 618 => 0, 619 => 0, 620 => 0, 621 => 0, 622 => 1, 623 => 0, 624 => 0, 625 => 0, 626 => 0, 627 => 0, 628 => 0, 629 => 0, 630 => 0, 631 => 1, 632 => 0, 633 => 0, 634 => 0, 635 => 0, 636 => 0, 637 => 0, 638 => 0, 639 => 0, 640 => 0, 641 => 0, 642 => 0, 643 => 0, 644 => 0, 645 => 0, 646 => 0, 647 => 0, 648 => 0, 649 => 0, 650 => 1, 651 => 0, 652 => 0, 653 => 0, 654 => 0, 655 => 0, 656 => 0, 657 => 0, 658 => 0, 659 => 1, 660 => 1, 661 => 1, 662 => 1, 663 => 1, 664 => 1, 665 => 1, 666 => 1, 667 => 1, 668 => 1, 669 => 0, 670 => 0, 671 => 0, 672 => 0, 673 => 0, 674 => 0, 675 
=> 1, 676 => 1, 677 => 1, 678 => 1, 679 => 1, 680 => 1, 681 => 1, 682 => 1, 683 => 1, 684 => 1, 685 => 1, 686 => 1, 687 => 1, 688 => 0, 689 => 0, 690 => 0, 691 => 0, 692 => 0, 693 => 0, 694 => 0, 695 => 0, 696 => 0, 697 => 1, 698 => 1, 699 => 1, 700 => 1, 701 => 1, 702 => 1, 703 => 1, 704 => 1, 705 => 1, 706 => 1, 707 => 0, 708 => 0, 709 => 0, 710 => 0, 711 => 0, 712 => 0, 713 => 0, 714 => 0, 715 => 0, 716 => 0, 717 => 0, 718 => 0, 719 => 0, 720 => 
0, 721 => 0, 722 => 1, 723 => 1, 724 => 1, 725 => 1, 726 => 1, 727 => 1, 728 => 1, 729 => 1, 730 => 1, 731 => 1, 732 => 1, 733 => 0, 734 => 0, 735 => 0, 736 => 0, 737 => 0, 738 => 0, 739 => 1, 740 => 1, 741 => 1, 742 => 0, 743 => 0, 744 => 0, 745 => 0, 746 => 0, 747 => 0, 748 => 1, 749 => 1, 750 => 1, 751 => 1, 752 => 1, 753 => 1, 754 => 1, 755 => 1, 756 => 1, 757 => 1, 758 => 0, 759 => 0, 760 => 0, 761 => 0, 762 => 0, 763 => 0, 764 => 0, 765 => 1, 
766 => 1, 767 => 1, 768 => 0, 769 => 0, 770 => 0, 771 => 0, 772 => 0, 773 => 0, 774 => 0, 775 => 0, 776 => 0, 777 => 1, 778 => 1, 779 => 1, 780 => 0, 781 => 0, 782 => 0, 783 => 0, 784 => 0, 785 => 0, 786 => 1, 787 => 1, 788 => 1, 789 => 1, 790 => 1, 791 => 1, 792 => 1, 793 => 1, 794 => 1, 795 => 1, 796 => 0, 797 => 0, 798 => 0, 799 => 0, 800 => 0, 801 => 0, 802 => 1, 803 => 1, 804 => 1, 805 => 1, 806 => 0, 807 => 0, 808 => 0, 809 => 1, 810 => 1, 811 => 1, 812 => 1, 813 => 1, 814 => 1, 815 => 0, 816 => 0, 817 => 0, 818 => 0, 819 => 0, 820 => 0, 821 => 0, 822 => 0, 823 => 1, 824 => 0, 825 => 0, 826 
=> 0, 827 => 0, 828 => 0, 829 => 0, 830 => 0, 831 => 0, 832 => 1, 833 => 0, 834 => 0, 835 => 0, 836 => 0, 837 => 0, 838 => 0, 839 => 1, 840 => 1, 841 => 1, 842 => 1, 843 => 0, 844 => 0, 845 => 0, 846 => 0, 847 => 0, 848 => 0, 849 => 0, 850 => 0, 851 => 1, 852 => 0, 853 => 0, 854 => 0, 855 => 0, 856 => 0, 857 => 0, 858 => 0, 859 => 0, 860 => 1, 861 => 0, 862 => 0, 863 => 0, 864 => 0, 865 => 0, 866 => 0, 867 => 0, 868 => 0, 869 => 0, 870 => 1, 871 => 
0, 872 => 0, 873 => 0, 874 => 0, 875 => 0, 876 => 0, 877 => 0, 878 => 0, 879 => 0, 880 => 0, 881 => 0, 882 => 0, 883 => 0, 884 => 0, 885 => 0, 886 => 1, 887 => 0, 888 => 0, 889 => 0, 890 => 0, 891 => 0, 892 => 0, 893 => 0, 894 => 0, 895 => 0, 896 => 1, 897 => 0, 898 => 0, 899 => 0, 900 => 0, 901 => 0, 902 => 0, 903 => 1, 904 => 1, 905 => 1, 906 => 0, 907 => 0, 908 => 0, 909 => 0, 910 => 0, 911 => 0, 912 => 0, 913 => 0, 914 => 0, 915 => 0, 916 => 0, 
917 => 0, 918 => 0, 919 => 0, 920 => 0, 921 => 0, 922 => 1, 923 => 0, 924 => 0, 925 => 0, 926 => 0, 927 => 0, 928 => 0, 929 => 1, 930 => 1, 931 => 1, 932 => 0, 933 => 0, 934 => 0, 935 => 0, 936 => 0, 937 => 0, 938 => 0, 939 => 0, 940 => 0, 941 => 1, 942 => 1, 943 => 1, 944 => 0, 945 => 0, 946 => 0, 947 => 0, 948 => 0, 949 => 0, 950 => 1, 951 => 0, 952 => 0, 953 => 0, 954 => 0, 955 => 0, 956 => 0, 957 => 0, 958 => 0, 959 => 1, 960 => 0, 961 => 0, 962 => 0, 963 => 0, 964 => 0, 965 => 0, 966 => 0, 967 => 0, 968 => 0, 969 => 1, 970 => 0, 971 => 0, 972 => 0, 973 => 0, 974 => 0, 975 => 0, 976 => 0, 977 
=> 0, 978 => 1, 979 => 0, 980 => 0, 981 => 0, 982 => 0, 983 => 0, 984 => 0, 985 => 1, 986 => 1, 987 => 1, 988 => 0, 989 => 0, 990 => 0, 991 => 0, 992 => 0, 993 => 0, 994 => 0, 995 => 0, 996 => 1, 997 => 1, 998 => 1, 999 => 1, 1000 => 0, 1001 => 0, 1002 => 0, 1003 => 1, 1004 => 1, 1005 => 1, 1006 => 0, 1007 => 0, 1008 => 0, 1009 => 0, 1010 => 0, 1011 => 0, 1012 => 0, 1013 => 0, 1014 => 0, 1015 => 1, 1016 => 1, 1017 => 1, 1018 => 0, 1019 => 0, 1020 => 0, 1021 => 0, 1022 => 1, 1023 => 1, 1024 => 1, 1025 => 0, 1026 => 0, 1027 => 0, 1028 => 0, 1029 => 0, 1030 => 0, 1031 => 0, 1032 => 0, 1033 => 0, 1034 => 1, 1035 => 1, 1036 => 1, 1037 => 0, 1038 => 0, 1039 => 0, 1040 => 0, 1041 => 0, 1042 => 0, 1043 => 0, 1044 => 0, 1045 => 0, 1046 => 0, 1047 => 0, 1048 => 1, 1049 => 1, 1050 => 1, 1051 => 0, 1052 => 0, 1053 => 0, 1054 => 0, 1055 => 0, 1056 => 0, 1057 => 0, 1058 => 0, 1059 => 0, 1060 => 1, 1061 => 1, 1062 => 1, 1063 => 0, 1064 => 0, 1065 => 0, 1066 => 0, 1067 => 1, 1068 => 1, 1069 => 1, 1070 => 0, 1071 => 0, 1072 => 0, 1073 => 0, 1074 => 0, 1075 => 0, 1076 => 0, 1077 => 0, 1078 => 0, 1079 => 0, 1080 => 0, 1081 => 0, 1082 => 0, 1083 => 0, 1084 => 0, 1085 => 0, 1086 => 1, 1087 => 1, 1088 => 1, 1089 => 0, 1090 => 0, 1091 => 0, 1092 => 0, 1093 => 1, 1094 => 1, 1095 => 1, 1096 => 0, 1097 => 0, 1098 => 0, 1099 => 0, 1100 => 0, 1101 => 0, 1102 => 0, 
1103 => 0, 1104 => 0, 1105 => 1, 1106 => 1, 1107 => 1, 1108 => 0, 1109 => 0, 1110 => 0, 1111 => 0, 1112 => 1, 1113 => 1, 1114 => 1, 1115 => 0, 1116 => 
0, 1117 => 0, 1118 => 0, 1119 => 0, 1120 => 0, 1121 => 0, 1122 => 0, 1123 => 1, 1124 => 1, 1125 => 1, 1126 => 1, 1127 => 0, 1128 => 0, 1129 => 0, 1130 
=> 0, 1131 => 0, 1132 => 0, 1133 => 1, 1134 => 1, 1135 => 1, 1136 => 0, 1137 => 0, 1138 => 0, 1139 => 0, 1140 => 0, 1141 => 0, 1142 => 1, 1143 => 1, 1144 => 1, 1145 => 0, 1146 => 0, 1147 => 0, 1148 => 0, 1149 => 1, 1150 => 1, 1151 => 1, 1152 => 0, 1153 => 0, 1154 => 0, 1155 => 0, 1156 => 0, 1157 => 0, 1158 => 0, 1159 => 0, 1160 => 1, 1161 => 1, 1162 => 1, 1163 => 0, 1164 => 0, 1165 => 0, 1166 => 0, 1167 => 1, 1168 => 1, 1169 => 1, 1170 => 0, 1171 => 0, 1172 => 0, 1173 => 0, 1174 => 0, 1175 => 0, 1176 => 0, 1177 => 0, 1178 => 0, 1179 => 1, 1180 => 1, 1181 => 1, 1182 => 0, 1183 => 0, 1184 => 0, 1185 => 0, 1186 => 1, 1187 => 1, 1188 => 1, 1189 => 0, 1190 => 0, 1191 => 0, 1192 => 0, 1193 => 0, 1194 => 0, 1195 => 0, 1196 => 0, 1197 => 0, 1198 => 1, 1199 => 1, 1200 => 1, 1201 => 0, 1202 => 0, 1203 => 0, 1204 => 0, 1205 => 0, 1206 => 0, 1207 => 0, 1208 => 0, 1209 => 0, 1210 => 0, 1211 => 0, 1212 => 1, 1213 => 1, 1214 => 1, 1215 => 0, 1216 => 0, 1217 => 0, 1218 => 0, 1219 => 0, 1220 => 0, 1221 => 0, 1222 => 0, 1223 => 0, 1224 => 1, 1225 => 1, 1226 => 1, 1227 => 0, 1228 => 0, 1229 => 0, 1230 => 0, 1231 => 1, 1232 => 1, 1233 => 1, 1234 => 0, 1235 => 0, 1236 => 0, 1237 => 0, 1238 => 0, 1239 => 0, 1240 => 0, 1241 => 0, 1242 => 0, 1243 => 0, 1244 => 0, 1245 => 0, 1246 => 0, 1247 => 0, 1248 => 0, 1249 => 0, 1250 => 1, 1251 => 1, 1252 => 1, 1253 => 0, 
1254 => 0, 1255 => 0, 1256 => 0, 1257 => 1, 1258 => 1, 1259 => 1, 1260 => 0, 1261 => 0, 1262 => 0, 1263 => 0, 1264 => 0, 1265 => 0, 1266 => 0, 1267 => 
0, 1268 => 0, 1269 => 1, 1270 => 1, 1271 => 1, 1272 => 0, 1273 => 0, 1274 => 0, 1275 => 0, 1276 => 1, 1277 => 1, 1278 => 1, 1279 => 0, 1280 => 0, 1281 
=> 0, 1282 => 0, 1283 => 0, 1284 => 0, 1285 => 0, 1286 => 0, 1287 => 1, 1288 => 1, 1289 => 1, 1290 => 0, 1291 => 0, 1292 => 0, 1293 => 0, 1294 => 0, 1295 => 0, 1296 => 0, 1297 => 1, 1298 => 1, 1299 => 1, 1300 => 0, 1301 => 0, 1302 => 0, 1303 => 0, 1304 => 0, 1305 => 0, 1306 => 1, 1307 => 1, 1308 => 1, 1309 => 0, 1310 => 0, 1311 => 0, 1312 => 0, 1313 => 1, 1314 => 1, 1315 => 1, 1316 => 0, 1317 => 0, 1318 => 0, 1319 => 0, 1320 => 0, 1321 => 0, 1322 => 0, 1323 => 0, 1324 => 1, 1325 => 1, 1326 => 1, 1327 => 0, 1328 => 0, 1329 => 0, 1330 => 0, 1331 => 1, 1332 => 1, 1333 => 1, 1334 => 0, 1335 => 0, 1336 => 0, 1337 => 0, 1338 => 0, 1339 => 0, 1340 => 0, 1341 => 0, 1342 => 0, 1343 => 1, 1344 => 1, 1345 => 1, 1346 => 0, 1347 => 0, 1348 => 0, 1349 => 0, 1350 => 1, 1351 => 1, 1352 => 1, 1353 => 0, 1354 => 0, 1355 => 0, 1356 => 0, 1357 => 0, 1358 => 0, 1359 => 0, 1360 => 0, 1361 => 0, 1362 => 1, 1363 => 1, 1364 => 1, 1365 => 0, 1366 => 0, 1367 => 0, 1368 => 0, 1369 => 0, 1370 => 0, 1371 => 0, 1372 => 0, 1373 => 0, 1374 => 0, 1375 => 0, 1376 => 1, 1377 => 1, 1378 => 1, 1379 => 0, 1380 => 0, 1381 => 0, 1382 => 0, 1383 => 0, 1384 => 0, 1385 => 0, 1386 => 0, 1387 => 0, 1388 => 1, 1389 => 1, 1390 => 1, 1391 => 0, 1392 => 0, 1393 => 0, 1394 => 0, 1395 => 1, 1396 => 1, 1397 => 1, 1398 => 0, 1399 => 0, 1400 => 0, 1401 => 0, 1402 => 0, 1403 => 0, 1404 => 1, 
1405 => 1, 1406 => 1, 1407 => 1, 1408 => 1, 1409 => 1, 1410 => 1, 1411 => 1, 1412 => 1, 1413 => 1, 1414 => 1, 1415 => 1, 1416 => 1, 1417 => 0, 1418 => 
0, 1419 => 0, 1420 => 0, 1421 => 1, 1422 => 1, 1423 => 1, 1424 => 0, 1425 => 0, 1426 => 0, 1427 => 0, 1428 => 0, 1429 => 0, 1430 => 0, 1431 => 0, 1432 
=> 0, 1433 => 1, 1434 => 1, 1435 => 1, 1436 => 0, 1437 => 0, 1438 => 0, 1439 => 0, 1440 => 1, 1441 => 1, 1442 => 1, 1443 => 0, 1444 => 0, 1445 => 0, 1446 => 0, 1447 => 0, 1448 => 0, 1449 => 0, 1450 => 0, 1451 => 1, 1452 => 1, 1453 => 1, 1454 => 0, 1455 => 0, 1456 => 0, 1457 => 0, 1458 => 0, 1459 => 0, 1460 => 0, 1461 => 1, 1462 => 1, 1463 => 1, 1464 => 0, 1465 => 0, 1466 => 0, 1467 => 0, 1468 => 0, 1469 => 0, 1470 => 1, 1471 => 1, 1472 => 1, 1473 => 0, 1474 => 0, 1475 => 0, 1476 => 0, 1477 => 1, 1478 => 1, 1479 => 1, 1480 => 0, 1481 => 0, 1482 => 0, 1483 => 0, 1484 => 0, 1485 => 0, 1486 => 0, 1487 => 0, 1488 => 1, 1489 => 1, 1490 => 1, 1491 => 0, 1492 => 0, 1493 => 0, 1494 => 0, 1495 => 1, 1496 => 1, 1497 => 1, 1498 => 0, 1499 => 0, 1500 => 0, 1501 => 0, 1502 => 0, 1503 => 0, 1504 => 0, 1505 => 0, 1506 => 0, 1507 => 1, 1508 => 1, 1509 => 1, 1510 => 0, 1511 => 0, 1512 => 0, 1513 => 0, 1514 => 1, 1515 => 1, 1516 => 1, 1517 => 0, 1518 => 0, 1519 => 0, 1520 => 0, 1521 => 0, 1522 => 0, 1523 => 0, 1524 => 0, 1525 => 0, 1526 => 1, 1527 => 1, 1528 => 1, 1529 => 0, 1530 => 0, 1531 => 0, 1532 => 0, 1533 => 0, 1534 => 0, 1535 => 0, 1536 => 0, 1537 => 0, 1538 => 0, 1539 => 0, 1540 => 1, 1541 => 1, 1542 => 1, 1543 => 0, 1544 => 0, 1545 => 0, 1546 => 0, 1547 => 0, 1548 => 0, 1549 => 0, 1550 => 0, 1551 => 0, 1552 => 1, 1553 => 1, 1554 => 1, 1555 => 0, 
1556 => 0, 1557 => 0, 1558 => 0, 1559 => 1, 1560 => 1, 1561 => 1, 1562 => 0, 1563 => 0, 1564 => 0, 1565 => 0, 1566 => 0, 1567 => 0, 1568 => 1, 1569 => 
1, 1570 => 1, 1571 => 1, 1572 => 1, 1573 => 1, 1574 => 1, 1575 => 1, 1576 => 1, 1577 => 1, 1578 => 1, 1579 => 1, 1580 => 1, 1581 => 0, 1582 => 0, 1583 
=> 0, 1584 => 0, 1585 => 1, 1586 => 1, 1587 => 1, 1588 => 0, 1589 => 0, 1590 => 0, 1591 => 0, 1592 => 0, 1593 => 0, 1594 => 0, 1595 => 0, 1596 => 0, 1597 => 1, 1598 => 1, 1599 => 1, 1600 => 0, 1601 => 0, 1602 => 0, 1603 => 0, 1604 => 1, 1605 => 1, 1606 => 1, 1607 => 0, 1608 => 0, 1609 => 0, 1610 => 0, 1611 => 0, 1612 => 0, 1613 => 0, 1614 => 0, 1615 => 1, 1616 => 1, 1617 => 1, 1618 => 1, 1619 => 0, 1620 => 0, 1621 => 0, 1622 => 0, 1623 => 0, 1624 => 0, 1625 => 1, 1626 => 1, 1627 => 1, 1628 => 0, 1629 => 0, 1630 => 0, 1631 => 0, 1632 => 0, 1633 => 0, 1634 => 1, 1635 => 1, 1636 => 1, 1637 => 0, 1638 => 0, 1639 => 0, 1640 => 0, 1641 => 1, 1642 => 1, 1643 => 1, 1644 => 0, 1645 => 0, 1646 => 0, 1647 => 0, 1648 => 0, 1649 => 0, 1650 => 0, 1651 => 0, 1652 => 1, 1653 => 1, 1654 => 1, 1655 => 0, 1656 => 0, 1657 => 0, 1658 => 0, 1659 => 1, 1660 => 1, 1661 => 1, 1662 => 0, 1663 => 0, 1664 => 0, 1665 => 0, 1666 => 0, 1667 => 0, 1668 => 0, 1669 => 0, 1670 => 0, 1671 => 1, 1672 => 1, 1673 => 1, 1674 => 0, 1675 => 0, 1676 => 0, 1677 => 0, 1678 => 1, 1679 => 1, 1680 => 1, 1681 => 1, 1682 => 0, 1683 => 0, 1684 => 0, 1685 => 0, 1686 => 0, 1687 => 0, 1688 => 0, 1689 => 1, 1690 => 1, 1691 => 0, 1692 => 0, 1693 => 0, 1694 => 0, 1695 => 0, 1696 => 0, 1697 => 0, 1698 => 0, 1699 => 0, 1700 => 0, 1701 => 0, 1702 => 0, 1703 => 0, 1704 => 1, 1705 => 1, 1706 => 1, 
1707 => 0, 1708 => 0, 1709 => 0, 1710 => 0, 1711 => 0, 1712 => 0, 1713 => 0, 1714 => 0, 1715 => 0, 1716 => 1, 1717 => 1, 1718 => 1, 1719 => 0, 1720 => 
0, 1721 => 0, 1722 => 0, 1723 => 1, 1724 => 1, 1725 => 1, 1726 => 0, 1727 => 0, 1728 => 0, 1729 => 0, 1730 => 0, 1731 => 0, 1732 => 1, 1733 => 0, 1734 
=> 0, 1735 => 0, 1736 => 0, 1737 => 0, 1738 => 0, 1739 => 0, 1740 => 0, 1741 => 0, 1742 => 1, 1743 => 1, 1744 => 1, 1745 => 0, 1746 => 0, 1747 => 0, 1748 => 0, 1749 => 0, 1750 => 0, 1751 => 1, 1752 => 0, 1753 => 0, 1754 => 0, 1755 => 0, 1756 => 0, 1757 => 0, 1758 => 0, 1759 => 0, 1760 => 1, 1761 => 1, 1762 => 1, 1763 => 1, 1764 => 0, 1765 => 0, 1766 => 0, 1767 => 0, 1768 => 1, 1769 => 1, 1770 => 1, 1771 => 0, 1772 => 0, 1773 => 0, 1774 => 0, 1775 => 0, 1776 => 0, 1777 => 0, 1778 => 0, 1779 => 1, 1780 => 0, 1781 => 0, 1782 => 0, 1783 => 0, 1784 => 0, 1785 => 0, 1786 => 0, 1787 => 0, 1788 => 0, 1789 => 1, 1790 => 1, 1791 => 1, 1792 => 0, 1793 => 0, 1794 => 0, 1795 => 0, 1796 => 0, 1797 => 0, 1798 => 0, 1799 => 0, 1800 => 0, 1801 => 0, 1802 => 0, 1803 => 0, 1804 => 0, 1805 => 1, 1806 => 1, 1807 => 1, 1808 => 0, 1809 => 0, 1810 => 0, 1811 => 0, 1812 => 0, 1813 => 0, 1814 => 0, 1815 => 0, 1816 => 1, 1817 => 1, 1818 => 1, 1819 => 0, 1820 => 0, 1821 => 0, 1822 => 0, 1823 => 1, 1824 => 1, 1825 => 1, 1826 => 0, 1827 => 0, 1828 => 0, 1829 => 0, 1830 => 0, 1831 => 0, 1832 => 0, 1833 => 0, 1834 => 0, 1835 => 1, 1836 => 1, 1837 => 1, 1838 => 0, 1839 => 0, 1840 => 0, 1841 => 0, 1842 => 1, 1843 => 1, 1844 => 1, 1845 => 1, 1846 => 1, 1847 => 1, 1848 => 1, 1849 => 1, 1850 => 1, 1851 => 1, 1852 => 1, 1853 => 1, 1854 => 1, 1855 => 0, 1856 => 0, 1857 => 0, 
1858 => 0, 1859 => 0, 1860 => 0, 1861 => 0, 1862 => 0, 1863 => 0, 1864 => 0, 1865 => 0, 1866 => 0, 1867 => 0, 1868 => 1, 1869 => 1, 1870 => 1, 1871 => 
0, 1872 => 0, 1873 => 0, 1874 => 0, 1875 => 0, 1876 => 0, 1877 => 0, 1878 => 0, 1879 => 0, 1880 => 1, 1881 => 1, 1882 => 1, 1883 => 0, 1884 => 0, 1885 
=> 0, 1886 => 0, 1887 => 1, 1888 => 1, 1889 => 1, 1890 => 0, 1891 => 0, 1892 => 0, 1893 => 0, 1894 => 1, 1895 => 1, 1896 => 1, 1897 => 0, 1898 => 0, 1899 => 0, 1900 => 0, 1901 => 0, 1902 => 0, 1903 => 0, 1904 => 0, 1905 => 0, 1906 => 1, 1907 => 1, 1908 => 1, 1909 => 0, 1910 => 0, 1911 => 0, 1912 => 0, 1913 => 0, 1914 => 0, 1915 => 1, 1916 => 1, 1917 => 1, 1918 => 1, 1919 => 1, 1920 => 1, 1921 => 1, 1922 => 1, 1923 => 1, 1924 => 1, 1925 => 1, 1926 => 1, 1927 => 1, 1928 => 0, 1929 => 0, 1930 => 0, 1931 => 0, 1932 => 1, 1933 => 1, 1934 => 1, 1935 => 1, 1936 => 1, 1937 => 1, 1938 => 1, 1939 => 1, 1940 => 1, 1941 => 1, 1942 => 1, 1943 => 1, 1944 => 0, 1945 => 0, 1946 => 0, 1947 => 0, 1948 => 0, 1949 => 0, 1950 => 0, 1951 => 0, 1952 => 0, 1953 => 1, 1954 => 1, 1955 => 1, 1956 => 0, 1957 => 0, 1958 => 0, 1959 => 0, 1960 => 0, 1961 => 0, 1962 => 0, 1963 => 0, 1964 => 0, 1965 => 0, 1966 => 0, 1967 => 0, 1968 => 0, 1969 => 1, 1970 => 1, 1971 => 1, 1972 => 0, 1973 => 0, 1974 => 0, 1975 => 0, 1976 => 0, 1977 => 0, 1978 => 0, 1979 => 0, 1980 => 1, 1981 => 1, 1982 => 1, 1983 => 0, 1984 => 0, 1985 => 0, 1986 => 0, 1987 => 1, 1988 => 1, 1989 => 1, 1990 => 0, 1991 => 0, 1992 => 0, 1993 => 0, 1994 => 0, 1995 => 0, 1996 => 0, 1997 => 0, 1998 => 0, 1999 => 1, 2000 => 1, 2001 => 1, 2002 => 0, 2003 => 0, 2004 => 0, 2005 => 0, 2006 => 1, 2007 => 1, 2008 => 1, 
2009 => 0, 2010 => 0, 2011 => 0, 2012 => 0, 2013 => 0, 2014 => 0, 2015 => 0, 2016 => 0, 2017 => 0, 2018 => 0, 2019 => 0, 2020 => 0, 2021 => 0, 2022 => 
0, 2023 => 0, 2024 => 0, 2025 => 0, 2026 => 0, 2027 => 0, 2028 => 0, 2029 => 0, 2030 => 0, 2031 => 0, 2032 => 1, 2033 => 1, 2034 => 1, 2035 => 0, 2036 
=> 0, 2037 => 0, 2038 => 0, 2039 => 0, 2040 => 0, 2041 => 0, 2042 => 0, 2043 => 0, 2044 => 1, 2045 => 0, 2046 => 0, 2047 => 0, 2048 => 0, 2049 => 0, 2050 => 0, 2051 => 1, 2052 => 1, 2053 => 1, 2054 => 0, 2055 => 0, 2056 => 0, 2057 => 0, 2058 => 1, 2059 => 1, 2060 => 1, 2061 => 0, 2062 => 0, 2063 => 0, 2064 => 0, 2065 => 0, 2066 => 0, 2067 => 0, 2068 => 0, 2069 => 0, 2070 => 1, 2071 => 1, 2072 => 1, 2073 => 0, 2074 => 0, 2075 => 0, 2076 => 0, 2077 => 0, 2078 => 0, 2079 => 0, 2080 => 0, 2081 => 0, 2082 => 0, 2083 => 0, 2084 => 0, 2085 => 0, 2086 => 0, 2087 => 0, 2088 => 1, 2089 => 1, 2090 => 1, 2091 => 1, 2092 => 0, 2093 => 0, 2094 => 0, 2095 => 0, 2096 => 1, 2097 => 1, 2098 => 1, 2099 => 0, 2100 => 0, 2101 => 0, 2102 => 0, 2103 => 0, 2104 => 0, 2105 => 0, 2106 => 0, 2107 => 0, 2108 => 0, 2109 => 0, 2110 => 0, 2111 => 0, 2112 => 0, 2113 => 0, 2114 => 0, 2115 => 0, 2116 => 0, 2117 => 1, 2118 => 1, 2119 => 1, 2120 => 0, 2121 => 0, 2122 => 0, 2123 => 0, 2124 => 0, 2125 => 0, 2126 => 0, 2127 => 0, 2128 => 0, 2129 => 0, 2130 => 0, 2131 => 0, 2132 => 0, 2133 => 1, 2134 => 1, 2135 => 1, 2136 => 0, 2137 => 0, 2138 => 0, 2139 => 0, 2140 => 0, 2141 => 0, 2142 => 0, 2143 => 0, 2144 => 1, 2145 => 1, 2146 => 1, 2147 => 0, 2148 => 0, 2149 => 0, 2150 => 0, 2151 => 1, 2152 => 1, 2153 => 1, 2154 => 0, 2155 => 0, 2156 => 0, 2157 => 0, 2158 => 0, 2159 => 0, 
2160 => 0, 2161 => 0, 2162 => 0, 2163 => 1, 2164 => 1, 2165 => 1, 2166 => 0, 2167 => 0, 2168 => 0, 2169 => 0, 2170 => 1, 2171 => 1, 2172 => 1, 2173 => 
0, 2174 => 0, 2175 => 0, 2176 => 0, 2177 => 0, 2178 => 0, 2179 => 0, 2180 => 0, 2181 => 0, 2182 => 0, 2183 => 0, 2184 => 0, 2185 => 0, 2186 => 0, 2187 
=> 0, 2188 => 0, 2189 => 0, 2190 => 0, 2191 => 0, 2192 => 0, 2193 => 0, 2194 => 0, 2195 => 0, 2196 => 1, 2197 => 1, 2198 => 1, 2199 => 1, 2200 => 1, 2201 => 1, 2202 => 1, 2203 => 1, 2204 => 1, 2205 => 1, 2206 => 1, 2207 => 1, 2208 => 1, 2209 => 0, 2210 => 0, 2211 => 0, 2212 => 0, 2213 => 0, 2214 => 0, 2215 => 1, 2216 => 1, 2217 => 1, 2218 => 0, 2219 => 0, 2220 => 0, 2221 => 0, 2222 => 1, 2223 => 1, 2224 => 1, 2225 => 0, 2226 => 0, 2227 => 0, 2228 => 0, 2229 => 0, 2230 => 0, 2231 => 0, 2232 => 0, 2233 => 0, 2234 => 1, 2235 => 1, 2236 => 1, 2237 => 0, 2238 => 0, 2239 => 0, 2240 => 0, 2241 => 0, 2242 => 0, 2243 => 0, 2244 => 0, 2245 => 0, 2246 => 0, 2247 => 0, 2248 => 0, 2249 => 0, 2250 => 0, 2251 => 0, 2252 => 0, 2253 => 1, 2254 => 1, 2255 => 1, 2256 => 0, 2257 => 0, 2258 => 0, 2259 => 0, 2260 => 1, 2261 => 1, 2262 => 1, 2263 => 0, 2264 => 0, 2265 => 0, 2266 => 0, 2267 => 0, 2268 => 0, 2269 => 0, 2270 => 0, 2271 => 0, 2272 => 0, 2273 => 0, 2274 => 0, 2275 => 0, 2276 => 0, 2277 => 0, 2278 => 0, 2279 => 0, 2280 => 0, 2281 => 1, 2282 => 1, 2283 => 1, 2284 => 0, 2285 => 0, 2286 => 0, 2287 => 0, 2288 => 0, 2289 => 0, 2290 => 0, 2291 => 0, 2292 => 0, 2293 => 0, 2294 => 0, 2295 => 0, 2296 => 0, 2297 => 0, 2298 => 1, 2299 => 1, 2300 => 0, 2301 => 0, 2302 => 0, 2303 => 0, 2304 => 0, 2305 => 0, 2306 => 0, 2307 => 0, 2308 => 1, 2309 => 1, 2310 => 0, 
2311 => 0, 2312 => 0, 2313 => 0, 2314 => 0, 2315 => 1, 2316 => 1, 2317 => 1, 2318 => 0, 2319 => 0, 2320 => 0, 2321 => 0, 2322 => 0, 2323 => 0, 2324 => 
0, 2325 => 0, 2326 => 0, 2327 => 1, 2328 => 1, 2329 => 1, 2330 => 0, 2331 => 0, 2332 => 0, 2333 => 0, 2334 => 1, 2335 => 0, 2336 => 1, 2337 => 0, 2338 
=> 0, 2339 => 0, 2340 => 0, 2341 => 0, 2342 => 0, 2343 => 0, 2344 => 0, 2345 => 0, 2346 => 0, 2347 => 0, 2348 => 0, 2349 => 0, 2350 => 0, 2351 => 0, 2352 => 0, 2353 => 0, 2354 => 0, 2355 => 0, 2356 => 0, 2357 => 0, 2358 => 0, 2359 => 0, 2360 => 1, 2361 => 1, 2362 => 1, 2363 => 1, 2364 => 0, 2365 => 0, 2366 => 0, 2367 => 0, 2368 => 0, 2369 => 0, 2370 => 0, 2371 => 0, 2372 => 0, 2373 => 0, 2374 => 0, 2375 => 0, 2376 => 0, 2377 => 0, 2378 => 0, 2379 => 1, 2380 => 1, 2381 => 1, 2382 => 0, 2383 => 0, 2384 => 0, 2385 => 0, 2386 => 1, 2387 => 1, 2388 => 1, 2389 => 0, 2390 => 0, 2391 => 0, 2392 => 0, 2393 => 0, 2394 => 0, 2395 => 0, 2396 => 0, 2397 => 0, 2398 => 0, 2399 => 1, 2400 => 1, 2401 => 0, 2402 => 0, 2403 => 0, 2404 => 0, 2405 => 0, 2406 => 0, 2407 => 0, 2408 => 0, 2409 => 0, 2410 => 0, 2411 => 0, 2412 => 0, 2413 => 0, 2414 => 0, 2415 => 0, 2416 => 0, 2417 => 1, 2418 => 0, 2419 => 1, 2420 => 0, 2421 => 0, 2422 => 0, 2423 => 0, 2424 => 0, 2425 => 1, 2426 => 1, 2427 => 0, 2428 => 0, 2429 => 0, 2430 => 0, 2431 => 0, 2432 => 0, 2433 => 0, 2434 => 0, 2435 => 0, 2436 => 0, 2437 => 0, 2438 => 0, 2439 => 0, 2440 => 0, 2441 => 0, 2442 => 0, 2443 => 0, 2444 => 0, 2445 => 1, 2446 => 1, 2447 => 1, 2448 => 0, 2449 => 0, 2450 => 0, 2451 => 0, 2452 => 0, 2453 => 0, 2454 => 0, 2455 => 0, 2456 => 0, 2457 => 0, 2458 => 0, 2459 => 0, 2460 => 0, 2461 => 0, 
2462 => 0, 2463 => 1, 2464 => 1, 2465 => 1, 2466 => 1, 2467 => 1, 2468 => 1, 2469 => 1, 2470 => 1, 2471 => 1, 2472 => 1, 2473 => 0, 2474 => 0, 2475 => 
0, 2476 => 0, 2477 => 0, 2478 => 0, 2479 => 1, 2480 => 1, 2481 => 1, 2482 => 0, 2483 => 0, 2484 => 0, 2485 => 0, 2486 => 0, 2487 => 0, 2488 => 0, 2489 
=> 0, 2490 => 0, 2491 => 1, 2492 => 1, 2493 => 1, 2494 => 0, 2495 => 0, 2496 => 0, 2497 => 0, 2498 => 0, 2499 => 0, 2500 => 0, 2501 => 1, 2502 => 1, 2503 => 1, 2504 => 1, 2505 => 1, 2506 => 1, 2507 => 1, 2508 => 1, 2509 => 1, 2510 => 1, 2511 => 0, 2512 => 0, 2513 => 0, 2514 => 0, 2515 => 0, 2516 => 0, 2517 => 0, 2518 => 0, 2519 => 0, 2520 => 0, 2521 => 0, 2522 => 0, 2523 => 0, 2524 => 1, 2525 => 1, 2526 => 1, 2527 => 0, 2528 => 0, 2529 => 0, 2530 => 0, 2531 => 0, 2532 => 0, 2533 => 0, 2534 => 0, 2535 => 0, 2536 => 0, 2537 => 0, 2538 => 0, 2539 => 0, 2540 => 0, 2541 => 0, 2542 => 0, 2543 => 1, 2544 => 1, 2545 => 1, 2546 => 0, 2547 => 0, 2548 => 0, 2549 => 0, 2550 => 0, 2551 => 0, 2552 => 1, 2553 => 1, 2554 => 1, 2555 => 1, 2556 => 1, 2557 => 1, 2558 => 1, 2559 => 1, 2560 => 0, 2561 => 0, 2562 => 0, 2563 => 0, 2564 => 1, 2565 => 0, 2566 => 0, 2567 => 0, 2568 => 0, 2569 => 0, 2570 => 0, 2571 => 1, 2572 => 1, 2573 => 1, 2574 => 1, 2575 => 1, 2576 => 1, 2577 => 1, 2578 => 1, 2579 => 1, 2580 => 1, 2581 => 0, 2582 => 0, 2583 => 0, 2584 => 0, 2585 => 0, 2586 => 0, 2587 => 0, 2588 => 0, 2589 => 0, 2590 => 1, 2591 => 1, 2592 => 1, 2593 => 1, 2594 => 1, 2595 => 1, 2596 => 1, 2597 => 1, 2598 => 1, 2599 => 1, 2600 => 0, 2601 => 0, 2602 => 0, 2603 => 0, 2604 => 0, 2605 => 0, 2606 => 0, 2607 => 0, 2608 => 0, 2609 => 1, 2610 => 1, 2611 => 1, 2612 => 0, 
2613 => 0, 2614 => 0, 2615 => 0, 2616 => 0, 2617 => 0, 2618 => 0, 2619 => 0, 2620 => 0, 2621 => 0, 2622 => 0, 2623 => 0, 2624 => 0, 2625 => 0, 2626 => 
0, 2627 => 1, 2628 => 1, 2629 => 1, 2630 => 1, 2631 => 1, 2632 => 1, 2633 => 1, 2634 => 1, 2635 => 1, 2636 => 1, 2637 => 0, 2638 => 0, 2639 => 0, 2640 
=> 0, 2641 => 0, 2642 => 0, 2643 => 1, 2644 => 1, 2645 => 1, 2646 => 1, 2647 => 0, 2648 => 0, 2649 => 0, 2650 => 0, 2651 => 0, 2652 => 0, 2653 => 0, 2654 => 0, 2655 => 1, 2656 => 1, 2657 => 1, 2658 => 0, 2659 => 0, 2660 => 0, 2661 => 0, 2662 => 0, 2663 => 0, 2664 => 1, 2665 => 1, 2666 => 1, 2667 => 1, 2668 => 1, 2669 => 1, 2670 => 1, 2671 => 1, 2672 => 1, 2673 => 1, 2674 => 1, 2675 => 0, 2676 => 0, 2677 => 0, 2678 => 0, 2679 => 0, 2680 => 0, 2681 => 0, 2682 => 0, 2683 => 0, 2684 => 0, 2685 => 0, 2686 => 0, 2687 => 0, 2688 => 1, 2689 => 1, 2690 => 1, 2691 => 0, 2692 => 0, 2693 => 0, 2694 => 0, 2695 => 0, 2696 => 0, 2697 => 0, 2698 => 0, 2699 => 0, 2700 => 0, 2701 => 0, 2702 => 0, 2703 => 0, 2704 => 0, 2705 => 0, 2706 => 0, 2707 => 1, 2708 => 1, 2709 => 1, 2710 => 0, 2711 => 0, 2712 => 0, 2713 => 0, 2714 => 0, 2715 => 0, 2716 => 1, 2717 => 1, 2718 => 1, 2719 => 1, 2720 => 1, 2721 => 1, 2722 => 1, 2723 => 1, 2724 => 0, 2725 => 0, 2726 => 0, 2727 => 0, 2728 => 1, 2729 => 0, 2730 => 0, 2731 => 0, 2732 => 0, 2733 => 0, 2734 => 0, 2735 => 1, 2736 => 1, 2737 => 1, 2738 => 1, 2739 => 1, 2740 => 1, 2741 => 1, 2742 => 1, 2743 => 1, 2744 => 1, 2745 => 0, 2746 => 0, 2747 => 0, 2748 => 0, 2749 => 0, 2750 => 0, 2751 => 0, 2752 => 0, 2753 => 0, 2754 => 1, 2755 => 1, 2756 => 1, 2757 => 1, 2758 => 1, 2759 => 1, 2760 => 1, 2761 => 1, 2762 => 1, 2763 => 1, 
2764 => 0, 2765 => 0, 2766 => 0, 2767 => 0, 2768 => 0, 2769 => 0, 2770 => 0, 2771 => 0, 2772 => 0, 2773 => 1, 2774 => 1, 2775 => 1, 2776 => 0, 2777 => 
0, 2778 => 0, 2779 => 0, 2780 => 0, 2781 => 0, 2782 => 0, 2783 => 0, 2784 => 0, 2785 => 0, 2786 => 0, 2787 => 0, 2788 => 0, 2789 => 0, 2790 => 0, 2791 
=> 0, 2792 => 0, 2793 => 0, 2794 => 0, 2795 => 0, 2796 => 0, 2797 => 0, 2798 => 0, 2799 => 0, 2800 => 0, 2801 => 0, 2802 => 0, 2803 => 0, 2804 => 0, 2805 => 0, 2806 => 0, 2807 => 0, 2808 => 0, 2809 => 0, 2810 => 0, 2811 => 0, 2812 => 0, 2813 => 0, 2814 => 0, 2815 => 0, 2816 => 0, 2817 => 0, 2818 => 0, 2819 => 0, 2820 => 0, 2821 => 0, 2822 => 0, 2823 => 0, 2824 => 0, 2825 => 0, 2826 => 0, 2827 => 0, 2828 => 0, 2829 => 0, 2830 => 0, 2831 => 0, 2832 => 0, 2833 => 0, 2834 => 0, 2835 => 0, 2836 => 0, 2837 => 0, 2838 => 0, 2839 => 0, 2840 => 0, 2841 => 0, 2842 => 0, 2843 => 0, 2844 => 0, 2845 => 0, 2846 => 0, 2847 => 0, 2848 => 0, 2849 => 0, 2850 => 0, 2851 => 0, 2852 => 0, 2853 => 0, 2854 => 0, 2855 => 0, 2856 => 0, 2857 => 0, 2858 => 0, 2859 => 0, 2860 => 0, 2861 => 0, 2862 => 0, 2863 => 0, 2864 => 0, 2865 => 0, 2866 => 0, 2867 => 0, 2868 => 0, 2869 => 0, 2870 => 0, 2871 => 0, 2872 => 0, 2873 => 0, 2874 => 0, 2875 => 0, 2876 => 0, 2877 => 0, 2878 => 0, 2879 => 0, 2880 => 0, 2881 => 0, 2882 => 0, 2883 => 0, 2884 => 0, 2885 => 0, 2886 => 0, 2887 => 0, 2888 => 0, 2889 => 0, 2890 => 0, 2891 => 0, 2892 => 0, 2893 => 0, 2894 => 0, 2895 => 0, 2896 => 0, 2897 => 0, 2898 => 0, 2899 => 0, 2900 => 0, 2901 => 0, 2902 => 0, 2903 => 0, 2904 => 0, 2905 => 0, 2906 => 0, 2907 => 0, 2908 => 0, 2909 => 0, 2910 => 0, 2911 => 0, 2912 => 0, 2913 => 0, 2914 => 0, 
2915 => 0, 2916 => 0, 2917 => 0, 2918 => 0, 2919 => 0, 2920 => 0, 2921 => 0, 2922 => 0, 2923 => 0, 2924 => 0, 2925 => 0, 2926 => 0, 2927 => 0, 2928 => 
0, 2929 => 0, 2930 => 0, 2931 => 0, 2932 => 0, 2933 => 0, 2934 => 0, 2935 => 0, 2936 => 0, 2937 => 0, 2938 => 0, 2939 => 0, 2940 => 0, 2941 => 0, 2942 
=> 0, 2943 => 0, 2944 => 0, 2945 => 0, 2946 => 0, 2947 => 0, 2948 => 0, 2949 => 0, 2950 => 0, 2951 => 0);

constant rom_option_2: rom_bitmap := (
0 => 0, 1 => 0, 2 => 0, 3 => 1, 4 => 1, 5 => 1, 6 => 0, 7 => 0, 8 => 0, 9 => 0, 10 => 0, 11 => 0, 12 => 0, 13 => 0, 14 => 0, 15 => 0, 16 => 0, 17 => 0, 18 => 0, 19 => 0, 20 => 0, 21 => 0, 22 => 0, 23 => 0, 24 => 0, 25 => 0, 26 => 0, 27 => 0, 28 => 0, 29 => 0, 30 => 0, 31 => 0, 32 => 0, 33 => 0, 34 => 
0, 35 => 0, 36 => 0, 37 => 0, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 0, 45 => 0, 46 => 0, 47 => 0, 48 => 0, 49 => 0, 50 => 0, 51 => 0, 52 => 0, 53 => 0, 54 => 0, 55 => 0, 56 => 0, 57 => 0, 58 => 0, 59 => 0, 60 => 0, 61 => 0, 62 => 0, 63 => 0, 64 => 0, 65 => 0, 66 => 0, 67 => 0, 68 => 0, 69 => 0, 70 => 0, 71 => 0, 72 => 0, 73 => 0, 74 => 0, 75 => 0, 76 => 0, 77 => 0, 78 => 0, 79 => 0, 80 => 0, 81 => 0, 82 => 0, 83 => 1, 84 => 1, 
85 => 1, 86 => 0, 87 => 0, 88 => 0, 89 => 0, 90 => 0, 91 => 0, 92 => 0, 93 => 0, 94 => 0, 95 => 0, 96 => 0, 97 => 0, 98 => 0, 99 => 0, 100 => 0, 101 => 0, 102 => 0, 103 => 0, 104 => 0, 105 => 0, 106 => 0, 107 => 0, 108 => 0, 109 => 0, 110 => 0, 111 => 0, 112 => 0, 113 => 0, 114 => 0, 115 => 0, 116 => 
0, 117 => 0, 118 => 0, 119 => 0, 120 => 0, 121 => 0, 122 => 0, 123 => 0, 124 => 0, 125 => 0, 126 => 0, 127 => 0, 128 => 0, 129 => 0, 130 => 0, 131 => 0, 132 => 0, 133 => 0, 134 => 0, 135 => 0, 136 => 0, 137 => 0, 138 => 0, 139 => 0, 140 => 0, 141 => 0, 142 => 0, 143 => 0, 144 => 0, 145 => 0, 146 => 0, 147 => 0, 148 => 0, 149 => 0, 150 => 0, 151 => 0, 152 => 0, 153 => 0, 154 => 0, 155 => 0, 156 => 0, 157 => 0, 158 => 0, 159 => 0, 160 => 0, 161 => 0, 
162 => 0, 163 => 0, 164 => 0, 165 => 0, 166 => 0, 167 => 1, 168 => 1, 169 => 1, 170 => 0, 171 => 0, 172 => 0, 173 => 0, 174 => 0, 175 => 0, 176 => 0, 177 => 0, 178 => 0, 179 => 0, 180 => 0, 181 => 0, 182 => 0, 183 => 0, 184 => 0, 185 => 0, 186 => 0, 187 => 0, 188 => 0, 189 => 0, 190 => 0, 191 => 0, 192 => 0, 193 => 0, 194 => 0, 195 => 0, 196 => 0, 197 => 0, 198 => 0, 199 => 0, 200 => 0, 201 => 0, 202 => 0, 203 => 0, 204 => 0, 205 => 0, 206 => 0, 207 => 0, 208 => 0, 209 => 0, 210 => 0, 211 => 0, 212 => 0, 213 => 0, 214 => 0, 215 => 0, 216 => 0, 217 => 0, 218 => 0, 219 => 0, 220 => 0, 221 => 0, 222 
=> 0, 223 => 0, 224 => 0, 225 => 0, 226 => 0, 227 => 0, 228 => 0, 229 => 0, 230 => 0, 231 => 0, 232 => 0, 233 => 0, 234 => 0, 235 => 0, 236 => 0, 237 => 0, 238 => 0, 239 => 0, 240 => 0, 241 => 0, 242 => 0, 243 => 0, 244 => 0, 245 => 0, 246 => 0, 247 => 1, 248 => 1, 249 => 1, 250 => 0, 251 => 0, 252 => 0, 253 => 0, 254 => 0, 255 => 0, 256 => 0, 257 => 0, 258 => 0, 259 => 0, 260 => 0, 261 => 0, 262 => 0, 263 => 0, 264 => 0, 265 => 0, 266 => 0, 267 => 
0, 268 => 0, 269 => 0, 270 => 0, 271 => 0, 272 => 0, 273 => 0, 274 => 0, 275 => 0, 276 => 0, 277 => 0, 278 => 0, 279 => 0, 280 => 0, 281 => 0, 282 => 0, 283 => 0, 284 => 0, 285 => 0, 286 => 0, 287 => 0, 288 => 0, 289 => 0, 290 => 0, 291 => 0, 292 => 0, 293 => 0, 294 => 0, 295 => 0, 296 => 0, 297 => 0, 298 => 0, 299 => 0, 300 => 0, 301 => 0, 302 => 0, 303 => 0, 304 => 0, 305 => 0, 306 => 0, 307 => 0, 308 => 0, 309 => 0, 310 => 0, 311 => 0, 312 => 0, 
313 => 0, 314 => 0, 315 => 0, 316 => 0, 317 => 0, 318 => 0, 319 => 0, 320 => 0, 321 => 0, 322 => 0, 323 => 0, 324 => 0, 325 => 0, 326 => 0, 327 => 0, 328 => 0, 329 => 0, 330 => 0, 331 => 1, 332 => 1, 333 => 1, 334 => 0, 335 => 0, 336 => 0, 337 => 0, 338 => 0, 339 => 0, 340 => 0, 341 => 0, 342 => 0, 343 => 0, 344 => 0, 345 => 0, 346 => 0, 347 => 0, 348 => 0, 349 => 0, 350 => 0, 351 => 0, 352 => 0, 353 => 0, 354 => 0, 355 => 0, 356 => 0, 357 => 0, 358 => 0, 359 => 0, 360 => 0, 361 => 0, 362 => 0, 363 => 0, 364 => 0, 365 => 0, 366 => 0, 367 => 0, 368 => 0, 369 => 0, 370 => 0, 371 => 0, 372 => 0, 373 
=> 0, 374 => 0, 375 => 0, 376 => 0, 377 => 0, 378 => 0, 379 => 0, 380 => 0, 381 => 0, 382 => 0, 383 => 0, 384 => 0, 385 => 0, 386 => 0, 387 => 0, 388 => 0, 389 => 0, 390 => 0, 391 => 0, 392 => 0, 393 => 0, 394 => 0, 395 => 0, 396 => 0, 397 => 0, 398 => 0, 399 => 0, 400 => 0, 401 => 0, 402 => 0, 403 => 0, 404 => 0, 405 => 0, 406 => 0, 407 => 0, 408 => 0, 409 => 0, 410 => 0, 411 => 1, 412 => 1, 413 => 1, 414 => 0, 415 => 0, 416 => 0, 417 => 0, 418 => 
0, 419 => 0, 420 => 0, 421 => 0, 422 => 0, 423 => 0, 424 => 0, 425 => 0, 426 => 0, 427 => 0, 428 => 0, 429 => 0, 430 => 0, 431 => 0, 432 => 0, 433 => 0, 434 => 0, 435 => 0, 436 => 0, 437 => 0, 438 => 0, 439 => 0, 440 => 0, 441 => 0, 442 => 0, 443 => 0, 444 => 0, 445 => 0, 446 => 0, 447 => 0, 448 => 0, 449 => 0, 450 => 0, 451 => 0, 452 => 0, 453 => 0, 454 => 0, 455 => 0, 456 => 0, 457 => 0, 458 => 0, 459 => 0, 460 => 0, 461 => 0, 462 => 0, 463 => 0, 
464 => 0, 465 => 0, 466 => 0, 467 => 0, 468 => 0, 469 => 0, 470 => 0, 471 => 0, 472 => 0, 473 => 0, 474 => 0, 475 => 0, 476 => 0, 477 => 0, 478 => 0, 479 => 0, 480 => 0, 481 => 0, 482 => 0, 483 => 0, 484 => 0, 485 => 0, 486 => 0, 487 => 0, 488 => 0, 489 => 0, 490 => 0, 491 => 0, 492 => 0, 493 => 0, 494 => 0, 495 => 1, 496 => 1, 497 => 1, 498 => 0, 499 => 0, 500 => 0, 501 => 0, 502 => 0, 503 => 0, 504 => 0, 505 => 0, 506 => 0, 507 => 0, 508 => 0, 509 => 0, 510 => 0, 511 => 1, 512 => 1, 513 => 1, 514 => 1, 515 => 0, 516 => 0, 517 => 0, 518 => 1, 519 => 0, 520 => 0, 521 => 0, 522 => 0, 523 => 1, 524 
=> 1, 525 => 1, 526 => 0, 527 => 0, 528 => 0, 529 => 0, 530 => 0, 531 => 0, 532 => 0, 533 => 1, 534 => 1, 535 => 1, 536 => 1, 537 => 1, 538 => 1, 539 => 1, 540 => 1, 541 => 1, 542 => 1, 543 => 0, 544 => 0, 545 => 0, 546 => 0, 547 => 0, 548 => 0, 549 => 0, 550 => 0, 551 => 0, 552 => 0, 553 => 0, 554 => 0, 555 => 0, 556 => 0, 557 => 0, 558 => 1, 559 => 1, 560 => 1, 561 => 1, 562 => 1, 563 => 1, 564 => 1, 565 => 1, 566 => 1, 567 => 1, 568 => 1, 569 => 
0, 570 => 0, 571 => 0, 572 => 0, 573 => 0, 574 => 0, 575 => 1, 576 => 1, 577 => 1, 578 => 0, 579 => 0, 580 => 0, 581 => 0, 582 => 0, 583 => 0, 584 => 1, 585 => 1, 586 => 1, 587 => 1, 588 => 1, 589 => 1, 590 => 1, 591 => 1, 592 => 1, 593 => 1, 594 => 1, 595 => 0, 596 => 0, 597 => 0, 598 => 0, 599 => 0, 600 => 0, 601 => 1, 602 => 1, 603 => 1, 604 => 0, 605 => 0, 606 => 0, 607 => 0, 608 => 0, 609 => 0, 610 => 0, 611 => 0, 612 => 1, 613 => 1, 614 => 1, 
615 => 1, 616 => 0, 617 => 0, 618 => 0, 619 => 0, 620 => 0, 621 => 0, 622 => 1, 623 => 1, 624 => 1, 625 => 1, 626 => 1, 627 => 1, 628 => 1, 629 => 1, 630 => 1, 631 => 1, 632 => 0, 633 => 0, 634 => 0, 635 => 0, 636 => 0, 637 => 0, 638 => 1, 639 => 1, 640 => 1, 641 => 1, 642 => 0, 643 => 0, 644 => 0, 645 => 1, 646 => 1, 647 => 1, 648 => 1, 649 => 1, 650 => 1, 651 => 0, 652 => 0, 653 => 0, 654 => 0, 655 => 0, 656 => 0, 657 => 0, 658 => 0, 659 => 1, 660 => 1, 661 => 1, 662 => 0, 663 => 0, 664 => 0, 665 => 0, 666 => 0, 667 => 0, 668 => 0, 669 => 0, 670 => 0, 671 => 0, 672 => 0, 673 => 0, 674 => 0, 675 
=> 1, 676 => 1, 677 => 1, 678 => 0, 679 => 0, 680 => 0, 681 => 0, 682 => 1, 683 => 0, 684 => 0, 685 => 0, 686 => 0, 687 => 1, 688 => 1, 689 => 1, 690 => 0, 691 => 0, 692 => 0, 693 => 0, 694 => 0, 695 => 0, 696 => 1, 697 => 1, 698 => 0, 699 => 0, 700 => 0, 701 => 0, 702 => 0, 703 => 0, 704 => 0, 705 => 0, 706 => 1, 707 => 0, 708 => 0, 709 => 0, 710 => 0, 711 => 0, 712 => 0, 713 => 0, 714 => 0, 715 => 0, 716 => 0, 717 => 0, 718 => 0, 719 => 0, 720 => 
0, 721 => 0, 722 => 1, 723 => 0, 724 => 0, 725 => 0, 726 => 0, 727 => 0, 728 => 0, 729 => 0, 730 => 0, 731 => 0, 732 => 1, 733 => 0, 734 => 0, 735 => 0, 736 => 0, 737 => 0, 738 => 0, 739 => 1, 740 => 1, 741 => 1, 742 => 0, 743 => 0, 744 => 0, 745 => 0, 746 => 0, 747 => 0, 748 => 0, 749 => 0, 750 => 0, 751 => 0, 752 => 0, 753 => 0, 754 => 0, 755 => 0, 756 => 0, 757 => 1, 758 => 0, 759 => 0, 760 => 0, 761 => 0, 762 => 0, 763 => 0, 764 => 0, 765 => 1, 
766 => 1, 767 => 1, 768 => 0, 769 => 0, 770 => 0, 771 => 0, 772 => 0, 773 => 0, 774 => 0, 775 => 0, 776 => 0, 777 => 1, 778 => 1, 779 => 1, 780 => 0, 781 => 0, 782 => 0, 783 => 0, 784 => 0, 785 => 0, 786 => 1, 787 => 0, 788 => 0, 789 => 0, 790 => 0, 791 => 0, 792 => 0, 793 => 0, 794 => 0, 795 => 1, 796 => 0, 797 => 0, 798 => 0, 799 => 0, 800 => 0, 801 => 0, 802 => 0, 803 => 0, 804 => 1, 805 => 1, 806 => 0, 807 => 0, 808 => 0, 809 => 0, 810 => 0, 811 => 0, 812 => 0, 813 => 0, 814 => 1, 815 => 0, 816 => 0, 817 => 0, 818 => 0, 819 => 0, 820 => 0, 821 => 1, 822 => 1, 823 => 1, 824 => 1, 825 => 1, 826 
=> 1, 827 => 1, 828 => 1, 829 => 1, 830 => 1, 831 => 1, 832 => 1, 833 => 1, 834 => 1, 835 => 1, 836 => 0, 837 => 0, 838 => 0, 839 => 1, 840 => 1, 841 => 1, 842 => 0, 843 => 0, 844 => 0, 845 => 0, 846 => 1, 847 => 0, 848 => 0, 849 => 0, 850 => 0, 851 => 1, 852 => 1, 853 => 1, 854 => 0, 855 => 0, 856 => 0, 857 => 0, 858 => 1, 859 => 1, 860 => 1, 861 => 0, 862 => 0, 863 => 0, 864 => 0, 865 => 0, 866 => 0, 867 => 0, 868 => 0, 869 => 0, 870 => 1, 871 => 
1, 872 => 1, 873 => 0, 874 => 0, 875 => 0, 876 => 0, 877 => 0, 878 => 0, 879 => 0, 880 => 0, 881 => 0, 882 => 0, 883 => 0, 884 => 1, 885 => 1, 886 => 1, 887 => 0, 888 => 0, 889 => 0, 890 => 0, 891 => 0, 892 => 0, 893 => 0, 894 => 0, 895 => 0, 896 => 1, 897 => 1, 898 => 1, 899 => 0, 900 => 0, 901 => 0, 902 => 0, 903 => 1, 904 => 1, 905 => 1, 906 => 0, 907 => 0, 908 => 0, 909 => 0, 910 => 0, 911 => 0, 912 => 0, 913 => 0, 914 => 0, 915 => 0, 916 => 0, 
917 => 0, 918 => 0, 919 => 0, 920 => 0, 921 => 0, 922 => 1, 923 => 1, 924 => 1, 925 => 0, 926 => 0, 927 => 0, 928 => 0, 929 => 1, 930 => 1, 931 => 1, 932 => 0, 933 => 0, 934 => 0, 935 => 0, 936 => 0, 937 => 0, 938 => 0, 939 => 0, 940 => 0, 941 => 1, 942 => 1, 943 => 1, 944 => 0, 945 => 0, 946 => 0, 947 => 0, 948 => 1, 949 => 1, 950 => 1, 951 => 0, 952 => 0, 953 => 0, 954 => 0, 955 => 0, 956 => 0, 957 => 0, 958 => 0, 959 => 1, 960 => 1, 961 => 1, 962 => 1, 963 => 0, 964 => 0, 965 => 0, 966 => 0, 967 => 0, 968 => 0, 969 => 1, 970 => 1, 971 => 1, 972 => 0, 973 => 0, 974 => 0, 975 => 0, 976 => 0, 977 
=> 0, 978 => 1, 979 => 1, 980 => 1, 981 => 0, 982 => 0, 983 => 0, 984 => 0, 985 => 1, 986 => 1, 987 => 1, 988 => 1, 989 => 1, 990 => 1, 991 => 1, 992 => 1, 993 => 1, 994 => 1, 995 => 1, 996 => 1, 997 => 1, 998 => 1, 999 => 1, 1000 => 0, 1001 => 0, 1002 => 0, 1003 => 1, 1004 => 1, 1005 => 1, 1006 => 0, 1007 => 0, 1008 => 0, 1009 => 0, 1010 => 1, 1011 => 0, 1012 => 0, 1013 => 0, 1014 => 0, 1015 => 1, 1016 => 1, 1017 => 1, 1018 => 0, 1019 => 0, 1020 => 0, 1021 => 0, 1022 => 1, 1023 => 1, 1024 => 1, 1025 => 0, 1026 => 0, 1027 => 0, 1028 => 0, 1029 => 0, 1030 => 0, 1031 => 0, 1032 => 0, 1033 => 0, 1034 => 1, 1035 => 1, 1036 => 1, 1037 => 0, 1038 => 0, 1039 => 0, 1040 => 0, 1041 => 0, 1042 => 0, 1043 => 0, 1044 => 0, 1045 => 0, 1046 => 0, 1047 => 0, 1048 => 1, 1049 => 1, 1050 => 1, 1051 => 0, 1052 => 0, 1053 => 0, 1054 => 0, 1055 => 0, 1056 => 0, 1057 => 0, 1058 => 0, 1059 => 0, 1060 => 1, 1061 => 1, 1062 => 1, 1063 => 0, 1064 => 0, 1065 => 0, 1066 => 0, 1067 => 1, 1068 => 1, 1069 => 1, 1070 => 0, 1071 => 0, 1072 => 0, 1073 => 0, 1074 => 0, 1075 => 0, 1076 => 0, 1077 => 0, 1078 => 0, 1079 => 0, 1080 => 0, 1081 => 0, 1082 => 0, 1083 => 0, 1084 => 0, 1085 => 0, 1086 => 1, 1087 => 1, 1088 => 1, 1089 => 0, 1090 => 0, 1091 => 0, 1092 => 0, 1093 => 1, 1094 => 1, 1095 => 1, 1096 => 0, 1097 => 0, 1098 => 0, 1099 => 0, 1100 => 0, 1101 => 0, 1102 => 0, 
1103 => 0, 1104 => 0, 1105 => 1, 1106 => 1, 1107 => 1, 1108 => 0, 1109 => 0, 1110 => 0, 1111 => 0, 1112 => 1, 1113 => 1, 1114 => 1, 1115 => 0, 1116 => 
0, 1117 => 0, 1118 => 0, 1119 => 0, 1120 => 0, 1121 => 0, 1122 => 0, 1123 => 1, 1124 => 1, 1125 => 1, 1126 => 0, 1127 => 0, 1128 => 0, 1129 => 0, 1130 
=> 0, 1131 => 0, 1132 => 0, 1133 => 1, 1134 => 1, 1135 => 1, 1136 => 0, 1137 => 0, 1138 => 0, 1139 => 0, 1140 => 0, 1141 => 0, 1142 => 1, 1143 => 1, 1144 => 1, 1145 => 0, 1146 => 0, 1147 => 0, 1148 => 0, 1149 => 0, 1150 => 0, 1151 => 1, 1152 => 1, 1153 => 1, 1154 => 0, 1155 => 0, 1156 => 0, 1157 => 0, 1158 => 0, 1159 => 0, 1160 => 0, 1161 => 0, 1162 => 0, 1163 => 0, 1164 => 0, 1165 => 0, 1166 => 0, 1167 => 1, 1168 => 1, 1169 => 1, 1170 => 0, 1171 => 0, 1172 => 0, 1173 => 0, 1174 => 1, 1175 => 0, 1176 => 0, 1177 => 0, 1178 => 0, 1179 => 1, 1180 => 1, 1181 => 1, 1182 => 0, 1183 => 0, 1184 => 0, 1185 => 0, 1186 => 1, 1187 => 1, 1188 => 1, 1189 => 0, 1190 => 0, 1191 => 0, 1192 => 0, 1193 => 0, 1194 => 0, 1195 => 0, 1196 => 0, 1197 => 0, 1198 => 1, 1199 => 1, 1200 => 1, 1201 => 0, 1202 => 0, 1203 => 0, 1204 => 0, 1205 => 0, 1206 => 0, 1207 => 0, 1208 => 0, 1209 => 0, 1210 => 0, 1211 => 0, 1212 => 1, 1213 => 1, 1214 => 1, 1215 => 0, 1216 => 0, 1217 => 0, 1218 => 0, 1219 => 0, 1220 => 0, 1221 => 0, 1222 => 0, 1223 => 0, 1224 => 1, 1225 => 1, 1226 => 1, 1227 => 0, 1228 => 0, 1229 => 0, 1230 => 0, 1231 => 1, 1232 => 1, 1233 => 1, 1234 => 0, 1235 => 0, 1236 => 0, 1237 => 0, 1238 => 0, 1239 => 0, 1240 => 1, 1241 => 1, 1242 => 1, 1243 => 1, 1244 => 1, 1245 => 1, 1246 => 1, 1247 => 1, 1248 => 1, 1249 => 1, 1250 => 1, 1251 => 1, 1252 => 1, 1253 => 0, 
1254 => 0, 1255 => 0, 1256 => 0, 1257 => 1, 1258 => 1, 1259 => 1, 1260 => 0, 1261 => 0, 1262 => 0, 1263 => 0, 1264 => 0, 1265 => 0, 1266 => 0, 1267 => 
0, 1268 => 0, 1269 => 1, 1270 => 1, 1271 => 1, 1272 => 0, 1273 => 0, 1274 => 0, 1275 => 0, 1276 => 1, 1277 => 1, 1278 => 1, 1279 => 0, 1280 => 0, 1281 
=> 0, 1282 => 0, 1283 => 0, 1284 => 0, 1285 => 0, 1286 => 0, 1287 => 1, 1288 => 1, 1289 => 1, 1290 => 0, 1291 => 0, 1292 => 0, 1293 => 0, 1294 => 0, 1295 => 0, 1296 => 0, 1297 => 1, 1298 => 1, 1299 => 1, 1300 => 0, 1301 => 0, 1302 => 0, 1303 => 0, 1304 => 0, 1305 => 0, 1306 => 1, 1307 => 1, 1308 => 1, 1309 => 0, 1310 => 0, 1311 => 0, 1312 => 0, 1313 => 0, 1314 => 0, 1315 => 1, 1316 => 1, 1317 => 1, 1318 => 0, 1319 => 0, 1320 => 0, 1321 => 0, 1322 => 0, 1323 => 0, 1324 => 0, 1325 => 0, 1326 => 0, 1327 => 0, 1328 => 0, 1329 => 0, 1330 => 0, 1331 => 1, 1332 => 1, 1333 => 1, 1334 => 0, 1335 => 0, 1336 => 0, 1337 => 0, 1338 => 1, 1339 => 0, 1340 => 0, 1341 => 0, 1342 => 0, 1343 => 1, 1344 => 1, 1345 => 1, 1346 => 0, 1347 => 0, 1348 => 0, 1349 => 0, 1350 => 1, 1351 => 1, 1352 => 1, 1353 => 0, 1354 => 0, 1355 => 0, 1356 => 0, 1357 => 0, 1358 => 0, 1359 => 0, 1360 => 0, 1361 => 0, 1362 => 1, 1363 => 1, 1364 => 1, 1365 => 0, 1366 => 0, 1367 => 0, 1368 => 0, 1369 => 0, 1370 => 0, 1371 => 0, 1372 => 0, 1373 => 0, 1374 => 0, 1375 => 0, 1376 => 1, 1377 => 1, 1378 => 1, 1379 => 0, 1380 => 0, 1381 => 0, 1382 => 0, 1383 => 0, 1384 => 0, 1385 => 0, 1386 => 0, 1387 => 0, 1388 => 1, 1389 => 1, 1390 => 1, 1391 => 0, 1392 => 0, 1393 => 0, 1394 => 0, 1395 => 1, 1396 => 1, 1397 => 1, 1398 => 0, 1399 => 0, 1400 => 0, 1401 => 0, 1402 => 0, 1403 => 0, 1404 => 1, 
1405 => 1, 1406 => 1, 1407 => 1, 1408 => 1, 1409 => 1, 1410 => 1, 1411 => 1, 1412 => 1, 1413 => 1, 1414 => 1, 1415 => 1, 1416 => 1, 1417 => 0, 1418 => 
0, 1419 => 0, 1420 => 0, 1421 => 1, 1422 => 1, 1423 => 1, 1424 => 0, 1425 => 0, 1426 => 0, 1427 => 0, 1428 => 0, 1429 => 0, 1430 => 0, 1431 => 0, 1432 
=> 0, 1433 => 1, 1434 => 1, 1435 => 1, 1436 => 0, 1437 => 0, 1438 => 0, 1439 => 0, 1440 => 1, 1441 => 1, 1442 => 1, 1443 => 0, 1444 => 0, 1445 => 0, 1446 => 0, 1447 => 0, 1448 => 0, 1449 => 0, 1450 => 0, 1451 => 1, 1452 => 1, 1453 => 1, 1454 => 1, 1455 => 0, 1456 => 0, 1457 => 0, 1458 => 0, 1459 => 0, 1460 => 0, 1461 => 1, 1462 => 1, 1463 => 1, 1464 => 0, 1465 => 0, 1466 => 0, 1467 => 0, 1468 => 0, 1469 => 0, 1470 => 1, 1471 => 1, 1472 => 1, 1473 => 0, 1474 => 0, 1475 => 0, 1476 => 0, 1477 => 0, 1478 => 0, 1479 => 1, 1480 => 1, 1481 => 1, 1482 => 0, 1483 => 0, 1484 => 0, 1485 => 0, 1486 => 0, 1487 => 0, 1488 => 0, 1489 => 0, 1490 => 0, 1491 => 0, 1492 => 0, 1493 => 0, 1494 => 0, 1495 => 1, 1496 => 1, 1497 => 1, 1498 => 0, 1499 => 0, 1500 => 0, 1501 => 0, 1502 => 1, 1503 => 0, 1504 => 0, 1505 => 0, 1506 => 0, 1507 => 1, 1508 => 1, 1509 => 1, 1510 => 0, 1511 => 0, 1512 => 0, 1513 => 0, 1514 => 1, 1515 => 1, 1516 => 1, 1517 => 0, 1518 => 0, 1519 => 0, 1520 => 0, 1521 => 0, 1522 => 0, 1523 => 0, 1524 => 0, 1525 => 0, 1526 => 1, 1527 => 1, 1528 => 1, 1529 => 0, 1530 => 0, 1531 => 0, 1532 => 0, 1533 => 0, 1534 => 0, 1535 => 0, 1536 => 0, 1537 => 0, 1538 => 0, 1539 => 0, 1540 => 1, 1541 => 1, 1542 => 1, 1543 => 0, 1544 => 0, 1545 => 0, 1546 => 0, 1547 => 0, 1548 => 0, 1549 => 0, 1550 => 0, 1551 => 0, 1552 => 1, 1553 => 1, 1554 => 1, 1555 => 0, 
1556 => 0, 1557 => 0, 1558 => 0, 1559 => 1, 1560 => 1, 1561 => 1, 1562 => 0, 1563 => 0, 1564 => 0, 1565 => 0, 1566 => 0, 1567 => 0, 1568 => 1, 1569 => 
0, 1570 => 0, 1571 => 0, 1572 => 0, 1573 => 0, 1574 => 0, 1575 => 0, 1576 => 0, 1577 => 0, 1578 => 1, 1579 => 1, 1580 => 1, 1581 => 0, 1582 => 0, 1583 
=> 0, 1584 => 0, 1585 => 0, 1586 => 0, 1587 => 1, 1588 => 0, 1589 => 0, 1590 => 0, 1591 => 0, 1592 => 0, 1593 => 0, 1594 => 0, 1595 => 0, 1596 => 1, 1597 => 1, 1598 => 1, 1599 => 1, 1600 => 0, 1601 => 0, 1602 => 0, 1603 => 0, 1604 => 1, 1605 => 1, 1606 => 1, 1607 => 0, 1608 => 0, 1609 => 0, 1610 => 0, 1611 => 0, 1612 => 0, 1613 => 0, 1614 => 0, 1615 => 1, 1616 => 0, 1617 => 0, 1618 => 0, 1619 => 0, 1620 => 0, 1621 => 0, 1622 => 0, 1623 => 0, 1624 => 0, 1625 => 1, 1626 => 1, 1627 => 1, 1628 => 0, 1629 => 0, 1630 => 0, 1631 => 0, 1632 => 0, 1633 => 0, 1634 => 0, 1635 => 0, 1636 => 0, 1637 => 0, 1638 => 0, 1639 => 0, 1640 => 0, 1641 => 0, 1642 => 0, 1643 => 1, 1644 => 1, 1645 => 1, 1646 => 0, 1647 => 0, 1648 => 0, 1649 => 0, 1650 => 0, 1651 => 0, 1652 => 1, 1653 => 1, 1654 => 1, 1655 => 1, 1656 => 0, 1657 => 0, 1658 => 0, 1659 => 1, 1660 => 1, 1661 => 1, 1662 => 0, 1663 => 0, 1664 => 0, 1665 => 0, 1666 => 1, 1667 => 0, 1668 => 0, 1669 => 0, 1670 => 0, 1671 => 1, 1672 => 1, 1673 => 1, 1674 => 0, 1675 => 0, 1676 => 0, 1677 => 0, 1678 => 1, 1679 => 1, 1680 => 1, 1681 => 0, 1682 => 0, 1683 => 0, 1684 => 0, 1685 => 0, 1686 => 0, 1687 => 0, 1688 => 0, 1689 => 0, 1690 => 1, 1691 => 1, 1692 => 1, 1693 => 0, 1694 => 0, 1695 => 0, 1696 => 0, 1697 => 0, 1698 => 0, 1699 => 0, 1700 => 0, 1701 => 0, 1702 => 0, 1703 => 0, 1704 => 1, 1705 => 1, 1706 => 1, 
1707 => 0, 1708 => 0, 1709 => 0, 1710 => 0, 1711 => 0, 1712 => 0, 1713 => 0, 1714 => 0, 1715 => 0, 1716 => 1, 1717 => 1, 1718 => 1, 1719 => 0, 1720 => 
0, 1721 => 0, 1722 => 0, 1723 => 1, 1724 => 1, 1725 => 1, 1726 => 0, 1727 => 0, 1728 => 0, 1729 => 0, 1730 => 1, 1731 => 1, 1732 => 1, 1733 => 0, 1734 
=> 0, 1735 => 0, 1736 => 0, 1737 => 0, 1738 => 0, 1739 => 0, 1740 => 0, 1741 => 0, 1742 => 1, 1743 => 1, 1744 => 1, 1745 => 0, 1746 => 0, 1747 => 0, 1748 => 0, 1749 => 0, 1750 => 0, 1751 => 1, 1752 => 1, 1753 => 1, 1754 => 1, 1755 => 1, 1756 => 1, 1757 => 1, 1758 => 1, 1759 => 1, 1760 => 1, 1761 => 1, 1762 => 1, 1763 => 1, 1764 => 0, 1765 => 0, 1766 => 0, 1767 => 0, 1768 => 1, 1769 => 1, 1770 => 1, 1771 => 1, 1772 => 1, 1773 => 1, 1774 => 1, 1775 => 1, 1776 => 1, 1777 => 1, 1778 => 1, 1779 => 1, 1780 => 0, 1781 => 0, 1782 => 0, 1783 => 0, 1784 => 0, 1785 => 0, 1786 => 0, 1787 => 0, 1788 => 0, 1789 => 1, 1790 => 1, 1791 => 1, 1792 => 0, 1793 => 0, 1794 => 0, 1795 => 0, 1796 => 0, 1797 => 0, 1798 => 0, 1799 => 0, 1800 => 0, 1801 => 0, 1802 => 0, 1803 => 0, 1804 => 0, 1805 => 0, 1806 => 0, 1807 => 1, 1808 => 1, 1809 => 1, 1810 => 0, 1811 => 0, 1812 => 0, 1813 => 0, 1814 => 0, 1815 => 0, 1816 => 1, 1817 => 1, 1818 => 1, 1819 => 0, 1820 => 0, 1821 => 0, 1822 => 0, 1823 => 1, 1824 => 1, 1825 => 1, 1826 => 0, 1827 => 0, 1828 => 0, 1829 => 0, 1830 => 1, 1831 => 0, 1832 => 0, 1833 => 0, 1834 => 0, 1835 => 1, 1836 => 1, 1837 => 1, 1838 => 0, 1839 => 0, 1840 => 0, 1841 => 0, 1842 => 1, 1843 => 1, 1844 => 1, 1845 => 0, 1846 => 0, 1847 => 0, 1848 => 0, 1849 => 0, 1850 => 0, 1851 => 0, 1852 => 0, 1853 => 0, 1854 => 1, 1855 => 1, 1856 => 1, 1857 => 0, 
1858 => 0, 1859 => 0, 1860 => 0, 1861 => 0, 1862 => 0, 1863 => 0, 1864 => 0, 1865 => 0, 1866 => 0, 1867 => 0, 1868 => 1, 1869 => 1, 1870 => 1, 1871 => 
0, 1872 => 0, 1873 => 0, 1874 => 0, 1875 => 0, 1876 => 0, 1877 => 0, 1878 => 0, 1879 => 0, 1880 => 1, 1881 => 0, 1882 => 0, 1883 => 0, 1884 => 0, 1885 
=> 0, 1886 => 0, 1887 => 1, 1888 => 1, 1889 => 1, 1890 => 0, 1891 => 0, 1892 => 0, 1893 => 0, 1894 => 1, 1895 => 1, 1896 => 1, 1897 => 0, 1898 => 0, 1899 => 0, 1900 => 0, 1901 => 0, 1902 => 0, 1903 => 0, 1904 => 0, 1905 => 0, 1906 => 1, 1907 => 1, 1908 => 1, 1909 => 0, 1910 => 0, 1911 => 0, 1912 => 0, 1913 => 0, 1914 => 0, 1915 => 0, 1916 => 0, 1917 => 0, 1918 => 0, 1919 => 0, 1920 => 0, 1921 => 0, 1922 => 0, 1923 => 0, 1924 => 1, 1925 => 1, 1926 => 1, 1927 => 1, 1928 => 0, 1929 => 0, 1930 => 0, 1931 => 0, 1932 => 1, 1933 => 1, 1934 => 1, 1935 => 0, 1936 => 0, 1937 => 0, 1938 => 0, 1939 => 0, 1940 => 0, 1941 => 0, 1942 => 0, 1943 => 0, 1944 => 0, 1945 => 0, 1946 => 0, 1947 => 0, 1948 => 0, 1949 => 0, 1950 => 0, 1951 => 0, 1952 => 0, 1953 => 1, 1954 => 1, 1955 => 1, 1956 => 0, 1957 => 0, 1958 => 0, 1959 => 0, 1960 => 0, 1961 => 0, 1962 => 0, 1963 => 0, 1964 => 0, 1965 => 0, 1966 => 0, 1967 => 0, 1968 => 0, 1969 => 0, 1970 => 0, 1971 => 1, 1972 => 1, 1973 => 1, 1974 => 0, 1975 => 0, 1976 => 0, 1977 => 0, 1978 => 0, 1979 => 0, 1980 => 1, 1981 => 1, 1982 => 1, 1983 => 0, 1984 => 0, 1985 => 0, 1986 => 0, 1987 => 1, 1988 => 1, 1989 => 1, 1990 => 0, 1991 => 0, 1992 => 0, 1993 => 0, 1994 => 1, 1995 => 0, 1996 => 0, 1997 => 0, 1998 => 0, 1999 => 1, 2000 => 1, 2001 => 1, 2002 => 0, 2003 => 0, 2004 => 0, 2005 => 0, 2006 => 1, 2007 => 1, 2008 => 1, 
2009 => 0, 2010 => 0, 2011 => 0, 2012 => 0, 2013 => 0, 2014 => 0, 2015 => 0, 2016 => 0, 2017 => 0, 2018 => 1, 2019 => 1, 2020 => 1, 2021 => 0, 2022 => 
0, 2023 => 0, 2024 => 0, 2025 => 0, 2026 => 0, 2027 => 0, 2028 => 0, 2029 => 0, 2030 => 0, 2031 => 0, 2032 => 1, 2033 => 1, 2034 => 1, 2035 => 1, 2036 
=> 1, 2037 => 1, 2038 => 1, 2039 => 1, 2040 => 1, 2041 => 1, 2042 => 1, 2043 => 1, 2044 => 1, 2045 => 0, 2046 => 0, 2047 => 0, 2048 => 0, 2049 => 0, 2050 => 0, 2051 => 1, 2052 => 1, 2053 => 1, 2054 => 0, 2055 => 0, 2056 => 0, 2057 => 0, 2058 => 1, 2059 => 1, 2060 => 1, 2061 => 0, 2062 => 0, 2063 => 0, 2064 => 0, 2065 => 0, 2066 => 0, 2067 => 0, 2068 => 0, 2069 => 0, 2070 => 1, 2071 => 1, 2072 => 1, 2073 => 0, 2074 => 0, 2075 => 0, 2076 => 0, 2077 => 0, 2078 => 0, 2079 => 0, 2080 => 0, 2081 => 0, 2082 => 0, 2083 => 0, 2084 => 0, 2085 => 0, 2086 => 0, 2087 => 0, 2088 => 0, 2089 => 1, 2090 => 1, 2091 => 1, 2092 => 0, 2093 => 0, 2094 => 0, 2095 => 0, 2096 => 1, 2097 => 1, 2098 => 1, 2099 => 0, 2100 => 0, 2101 => 0, 2102 => 0, 2103 => 0, 2104 => 0, 2105 => 0, 2106 => 0, 2107 => 0, 2108 => 0, 2109 => 0, 2110 => 0, 2111 => 0, 2112 => 0, 2113 => 0, 2114 => 0, 2115 => 0, 2116 => 0, 2117 => 1, 2118 => 1, 2119 => 1, 2120 => 0, 2121 => 0, 2122 => 0, 2123 => 0, 2124 => 0, 2125 => 0, 2126 => 0, 2127 => 0, 2128 => 0, 2129 => 0, 2130 => 0, 2131 => 0, 2132 => 0, 2133 => 0, 2134 => 0, 2135 => 1, 2136 => 1, 2137 => 1, 2138 => 0, 2139 => 0, 2140 => 0, 2141 => 0, 2142 => 0, 2143 => 0, 2144 => 1, 2145 => 1, 2146 => 1, 2147 => 1, 2148 => 0, 2149 => 0, 2150 => 0, 2151 => 1, 2152 => 1, 2153 => 1, 2154 => 0, 2155 => 0, 2156 => 0, 2157 => 0, 2158 => 0, 2159 => 0, 
2160 => 0, 2161 => 0, 2162 => 0, 2163 => 1, 2164 => 1, 2165 => 1, 2166 => 0, 2167 => 0, 2168 => 0, 2169 => 0, 2170 => 1, 2171 => 1, 2172 => 1, 2173 => 
0, 2174 => 0, 2175 => 0, 2176 => 0, 2177 => 0, 2178 => 0, 2179 => 0, 2180 => 0, 2181 => 0, 2182 => 1, 2183 => 1, 2184 => 1, 2185 => 0, 2186 => 0, 2187 
=> 0, 2188 => 0, 2189 => 0, 2190 => 0, 2191 => 0, 2192 => 0, 2193 => 0, 2194 => 0, 2195 => 0, 2196 => 1, 2197 => 1, 2198 => 1, 2199 => 1, 2200 => 1, 2201 => 1, 2202 => 1, 2203 => 1, 2204 => 1, 2205 => 1, 2206 => 1, 2207 => 1, 2208 => 1, 2209 => 0, 2210 => 0, 2211 => 0, 2212 => 0, 2213 => 0, 2214 => 0, 2215 => 1, 2216 => 1, 2217 => 1, 2218 => 0, 2219 => 0, 2220 => 0, 2221 => 0, 2222 => 1, 2223 => 1, 2224 => 1, 2225 => 0, 2226 => 0, 2227 => 0, 2228 => 0, 2229 => 0, 2230 => 0, 2231 => 0, 2232 => 0, 2233 => 0, 2234 => 1, 2235 => 1, 2236 => 1, 2237 => 0, 2238 => 0, 2239 => 0, 2240 => 0, 2241 => 0, 2242 => 0, 2243 => 0, 2244 => 0, 2245 => 0, 2246 => 0, 2247 => 0, 2248 => 0, 2249 => 0, 2250 => 0, 2251 => 0, 2252 => 0, 2253 => 1, 2254 => 1, 2255 => 1, 2256 => 0, 2257 => 0, 2258 => 0, 2259 => 0, 2260 => 1, 2261 => 1, 2262 => 1, 2263 => 0, 2264 => 0, 2265 => 0, 2266 => 0, 2267 => 0, 2268 => 0, 2269 => 0, 2270 => 0, 2271 => 0, 2272 => 0, 2273 => 0, 2274 => 0, 2275 => 0, 2276 => 0, 2277 => 0, 2278 => 0, 2279 => 0, 2280 => 0, 2281 => 1, 2282 => 1, 2283 => 1, 2284 => 0, 2285 => 0, 2286 => 0, 2287 => 0, 2288 => 0, 2289 => 0, 2290 => 0, 2291 => 0, 2292 => 0, 2293 => 0, 2294 => 0, 2295 => 0, 2296 => 0, 2297 => 0, 2298 => 0, 2299 => 0, 2300 => 0, 2301 => 1, 2302 => 1, 2303 => 1, 2304 => 1, 2305 => 1, 2306 => 1, 2307 => 1, 2308 => 1, 2309 => 0, 2310 => 0, 
2311 => 0, 2312 => 0, 2313 => 0, 2314 => 0, 2315 => 0, 2316 => 0, 2317 => 0, 2318 => 1, 2319 => 1, 2320 => 1, 2321 => 1, 2322 => 1, 2323 => 1, 2324 => 
1, 2325 => 1, 2326 => 1, 2327 => 1, 2328 => 0, 2329 => 0, 2330 => 0, 2331 => 0, 2332 => 0, 2333 => 0, 2334 => 0, 2335 => 0, 2336 => 0, 2337 => 1, 2338 
=> 1, 2339 => 1, 2340 => 1, 2341 => 1, 2342 => 1, 2343 => 1, 2344 => 1, 2345 => 1, 2346 => 1, 2347 => 0, 2348 => 0, 2349 => 0, 2350 => 0, 2351 => 0, 2352 => 0, 2353 => 0, 2354 => 0, 2355 => 0, 2356 => 0, 2357 => 0, 2358 => 0, 2359 => 0, 2360 => 1, 2361 => 1, 2362 => 1, 2363 => 0, 2364 => 0, 2365 => 0, 2366 => 0, 2367 => 0, 2368 => 0, 2369 => 0, 2370 => 0, 2371 => 0, 2372 => 0, 2373 => 0, 2374 => 0, 2375 => 0, 2376 => 0, 2377 => 0, 2378 => 0, 2379 => 1, 2380 => 1, 2381 => 1, 2382 => 0, 2383 => 0, 2384 => 0, 2385 => 0, 2386 => 0, 2387 => 0, 2388 => 1, 2389 => 1, 2390 => 1, 2391 => 1, 2392 => 1, 2393 => 1, 2394 => 1, 2395 => 1, 2396 => 0, 2397 => 0, 2398 => 0, 2399 => 0, 2400 => 1, 2401 => 0, 2402 => 0, 2403 => 0, 2404 => 0, 2405 => 0, 2406 => 0, 2407 => 1, 2408 => 1, 2409 => 1, 2410 => 1, 2411 => 1, 2412 => 1, 2413 => 1, 2414 => 1, 2415 => 1, 2416 => 1, 2417 => 0, 2418 => 0, 2419 => 0, 2420 => 0, 2421 => 0, 2422 => 0, 2423 => 0, 2424 => 0, 2425 => 0, 2426 => 1, 2427 => 1, 2428 => 1, 2429 => 1, 2430 => 1, 2431 => 1, 2432 => 1, 2433 => 1, 2434 => 1, 2435 => 1, 2436 => 0, 2437 => 0, 2438 => 0, 2439 => 0, 2440 => 0, 2441 => 0, 2442 => 0, 2443 => 0, 2444 => 0, 2445 => 1, 2446 => 1, 2447 => 1, 2448 => 0, 2449 => 0, 2450 => 0, 2451 => 0, 2452 => 0, 2453 => 0, 2454 => 0, 2455 => 0, 2456 => 0, 2457 => 0, 2458 => 0, 2459 => 0, 2460 => 0, 2461 => 0, 
2462 => 0, 2463 => 0, 2464 => 0, 2465 => 1, 2466 => 1, 2467 => 1, 2468 => 1, 2469 => 1, 2470 => 1, 2471 => 1, 2472 => 1, 2473 => 0, 2474 => 0, 2475 => 
0, 2476 => 0, 2477 => 0, 2478 => 0, 2479 => 0, 2480 => 0, 2481 => 0, 2482 => 1, 2483 => 1, 2484 => 1, 2485 => 1, 2486 => 1, 2487 => 1, 2488 => 1, 2489 
=> 1, 2490 => 1, 2491 => 1, 2492 => 0, 2493 => 0, 2494 => 0, 2495 => 0, 2496 => 0, 2497 => 0, 2498 => 0, 2499 => 0, 2500 => 1, 2501 => 1, 2502 => 1, 2503 => 1, 2504 => 1, 2505 => 1, 2506 => 1, 2507 => 1, 2508 => 1, 2509 => 1, 2510 => 1, 2511 => 0, 2512 => 0, 2513 => 0, 2514 => 0, 2515 => 0, 2516 => 0, 2517 => 0, 2518 => 0, 2519 => 0, 2520 => 0, 2521 => 0, 2522 => 0, 2523 => 0, 2524 => 1, 2525 => 1, 2526 => 1, 2527 => 0, 2528 => 0, 2529 => 0, 2530 => 0, 2531 => 0, 2532 => 0, 2533 => 0, 2534 => 0, 2535 => 0, 2536 => 0, 2537 => 0, 2538 => 0, 2539 => 0, 2540 => 0, 2541 => 0, 2542 => 0, 2543 => 1, 2544 => 1, 2545 => 1, 2546 => 0, 2547 => 0, 2548 => 0, 2549 => 0, 2550 => 0, 2551 => 0, 2552 => 1, 2553 => 1, 2554 => 1, 2555 => 1, 2556 => 1, 2557 => 1, 2558 => 1, 2559 => 1, 2560 => 0, 2561 => 0, 2562 => 0, 2563 => 0, 2564 => 1, 2565 => 0, 2566 => 0, 2567 => 0, 2568 => 0, 2569 => 0, 2570 => 0, 2571 => 1, 2572 => 1, 2573 => 1, 2574 => 1, 2575 => 1, 2576 => 1, 2577 => 1, 2578 => 1, 2579 => 1, 2580 => 1, 2581 => 0, 2582 => 0, 2583 => 0, 2584 => 0, 2585 => 0, 2586 => 0, 2587 => 0, 2588 => 0, 2589 => 0, 2590 => 1, 2591 => 1, 2592 => 1, 2593 => 1, 2594 => 1, 2595 => 1, 2596 => 1, 2597 => 1, 2598 => 1, 2599 => 1, 2600 => 0, 2601 => 0, 2602 => 0, 2603 => 0, 2604 => 0, 2605 => 0, 2606 => 0, 2607 => 0, 2608 => 0, 2609 => 1, 2610 => 1, 2611 => 1, 2612 => 0, 
2613 => 0, 2614 => 0, 2615 => 0, 2616 => 0, 2617 => 0, 2618 => 0, 2619 => 0, 2620 => 0, 2621 => 0, 2622 => 0, 2623 => 0, 2624 => 0, 2625 => 0, 2626 => 
0, 2627 => 0, 2628 => 0, 2629 => 0, 2630 => 0, 2631 => 0, 2632 => 0, 2633 => 0, 2634 => 0, 2635 => 0, 2636 => 0, 2637 => 0, 2638 => 0, 2639 => 0, 2640 
=> 0, 2641 => 0, 2642 => 0, 2643 => 0, 2644 => 0, 2645 => 0, 2646 => 0, 2647 => 0, 2648 => 0, 2649 => 0, 2650 => 0, 2651 => 0, 2652 => 0, 2653 => 0, 2654 => 0, 2655 => 0, 2656 => 0, 2657 => 0, 2658 => 0, 2659 => 0, 2660 => 0, 2661 => 0, 2662 => 0, 2663 => 0, 2664 => 0, 2665 => 0, 2666 => 0, 2667 => 0, 2668 => 0, 2669 => 0, 2670 => 0, 2671 => 0, 2672 => 0, 2673 => 0, 2674 => 0, 2675 => 0, 2676 => 0, 2677 => 0, 2678 => 0, 2679 => 0, 2680 => 0, 2681 => 0, 2682 => 0, 2683 => 0, 2684 => 0, 2685 => 0, 2686 => 0, 2687 => 0, 2688 => 0, 2689 => 0, 2690 => 0, 2691 => 0, 2692 => 0, 2693 => 0, 2694 => 0, 2695 => 0, 2696 => 0, 2697 => 0, 2698 => 0, 2699 => 0, 2700 => 0, 2701 => 0, 2702 => 0, 2703 => 0, 2704 => 0, 2705 => 0, 2706 => 0, 2707 => 0, 2708 => 0, 2709 => 0, 2710 => 0, 2711 => 0, 2712 => 0, 2713 => 0, 2714 => 0, 2715 => 0, 2716 => 0, 2717 => 0, 2718 => 0, 2719 => 0, 2720 => 0, 2721 => 0, 2722 => 0, 2723 => 0, 2724 => 0, 2725 => 0, 2726 => 0, 2727 => 0, 2728 => 0, 2729 => 0, 2730 => 0, 2731 => 0, 2732 => 0, 2733 => 0, 2734 => 0, 2735 => 0, 2736 => 0, 2737 => 0, 2738 => 0, 2739 => 0, 2740 => 0, 2741 => 0, 2742 => 0, 2743 => 0, 2744 => 0, 2745 => 0, 2746 => 0, 2747 => 0, 2748 => 0, 2749 => 0, 2750 => 0, 2751 => 0, 2752 => 0, 2753 => 0, 2754 => 0, 2755 => 0, 2756 => 0, 2757 => 0, 2758 => 0, 2759 => 0, 2760 => 0, 2761 => 0, 2762 => 0, 2763 => 0, 
2764 => 0, 2765 => 0, 2766 => 0, 2767 => 0, 2768 => 0, 2769 => 0, 2770 => 0, 2771 => 0, 2772 => 0, 2773 => 0, 2774 => 0, 2775 => 0, 2776 => 0, 2777 => 
0, 2778 => 0, 2779 => 0, 2780 => 0, 2781 => 0, 2782 => 0, 2783 => 0, 2784 => 0, 2785 => 0, 2786 => 0, 2787 => 0, 2788 => 0, 2789 => 0, 2790 => 0, 2791 
=> 0, 2792 => 0, 2793 => 0, 2794 => 0, 2795 => 0, 2796 => 0, 2797 => 0, 2798 => 0, 2799 => 0, 2800 => 0, 2801 => 0, 2802 => 0, 2803 => 0, 2804 => 0, 2805 => 0, 2806 => 0, 2807 => 0, 2808 => 0, 2809 => 0, 2810 => 0, 2811 => 0, 2812 => 0, 2813 => 0, 2814 => 0, 2815 => 0, 2816 => 0, 2817 => 0, 2818 => 0, 2819 => 0, 2820 => 0, 2821 => 0, 2822 => 0, 2823 => 0, 2824 => 0, 2825 => 0, 2826 => 0, 2827 => 0, 2828 => 0, 2829 => 0, 2830 => 0, 2831 => 0, 2832 => 0, 2833 => 0, 2834 => 0, 2835 => 0, 2836 => 0, 2837 => 0, 2838 => 0, 2839 => 0, 2840 => 0, 2841 => 0, 2842 => 0, 2843 => 0, 2844 => 0, 2845 => 0, 2846 => 0, 2847 => 0, 2848 => 0, 2849 => 0, 2850 => 0, 2851 => 0, 2852 => 0, 2853 => 0, 2854 => 0, 2855 => 0, 2856 => 0, 2857 => 0, 2858 => 0, 2859 => 0, 2860 => 0, 2861 => 0, 2862 => 0, 2863 => 0, 2864 => 0, 2865 => 0, 2866 => 0, 2867 => 0, 2868 => 0, 2869 => 0, 2870 => 0, 2871 => 0, 2872 => 0, 2873 => 0, 2874 => 0, 2875 => 0, 2876 => 0, 2877 => 0, 2878 => 0, 2879 => 0, 2880 => 0, 2881 => 0, 2882 => 0, 2883 => 0, 2884 => 0, 2885 => 0, 2886 => 0, 2887 => 0, 2888 => 0, 2889 => 0, 2890 => 0, 2891 => 0, 2892 => 0, 2893 => 0, 2894 => 0, 2895 => 0, 2896 => 0, 2897 => 0, 2898 => 0, 2899 => 0, 2900 => 0, 2901 => 0, 2902 => 0, 2903 => 0, 2904 => 0, 2905 => 0, 2906 => 0, 2907 => 0, 2908 => 0, 2909 => 0, 2910 => 0, 2911 => 0, 2912 => 0, 2913 => 0, 2914 => 0, 
2915 => 0, 2916 => 0, 2917 => 0, 2918 => 0, 2919 => 0, 2920 => 0, 2921 => 0, 2922 => 0, 2923 => 0, 2924 => 0, 2925 => 0, 2926 => 0, 2927 => 0, 2928 => 
0, 2929 => 0, 2930 => 0, 2931 => 0, 2932 => 0, 2933 => 0, 2934 => 0, 2935 => 0, 2936 => 0, 2937 => 0, 2938 => 0, 2939 => 0, 2940 => 0, 2941 => 0, 2942 
=> 0, 2943 => 0, 2944 => 0, 2945 => 0, 2946 => 0, 2947 => 0, 2948 => 0, 2949 => 0, 2950 => 0, 2951 => 0
);

constant rom_arrow: rom_bitmap_arrow := (

0 => 0, 1 => 0, 2 => 0, 3 => 0, 4 => 0, 5 => 0, 6 => 0, 7 => 0, 8 => 0, 9 => 0, 10 => 0, 11 => 0, 12 => 0, 13 => 0, 14 => 0, 15 => 0, 16 => 0, 17 => 0, 18 => 0, 19 => 0, 20 => 0, 21 => 0, 22 => 0, 23 => 0, 24 => 0, 25 => 0, 26 => 0, 27 => 0, 28 => 0, 29 => 0, 30 => 0, 31 => 0, 32 => 0, 33 => 0, 34 => 
0, 35 => 0, 36 => 0, 37 => 0, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 0, 45 => 0, 46 => 0, 47 => 0, 48 => 0, 49 => 0, 50 => 0, 51 => 1, 52 => 1, 53 => 1, 54 => 1, 55 => 0, 56 => 0, 57 => 0, 58 => 0, 59 => 0, 60 => 0, 61 => 0, 62 => 0, 63 => 0, 64 => 0, 65 => 0, 66 => 0, 67 => 0, 68 => 0, 69 => 0, 70 => 0, 71 => 0, 72 => 0, 73 => 0, 74 => 0, 75 => 0, 76 => 0, 77 => 0, 78 => 0, 79 => 0, 80 => 0, 81 => 0, 82 => 0, 83 => 0, 84 => 0, 
85 => 0, 86 => 0, 87 => 1, 88 => 1, 89 => 1, 90 => 1, 91 => 0, 92 => 0, 93 => 0, 94 => 0, 95 => 0, 96 => 0, 97 => 0, 98 => 0, 99 => 0, 100 => 0, 101 => 0, 102 => 0, 103 => 0, 104 => 0, 105 => 0, 106 => 0, 107 => 0, 108 => 0, 109 => 0, 110 => 0, 111 => 0, 112 => 0, 113 => 0, 114 => 0, 115 => 0, 116 => 
0, 117 => 0, 118 => 0, 119 => 0, 120 => 0, 121 => 1, 122 => 1, 123 => 1, 124 => 0, 125 => 0, 126 => 0, 127 => 0, 128 => 0, 129 => 0, 130 => 0, 131 => 0, 132 => 0, 133 => 0, 134 => 0, 135 => 0, 136 => 0, 137 => 0, 138 => 0, 139 => 0, 140 => 0, 141 => 0, 142 => 0, 143 => 0, 144 => 0, 145 => 0, 146 => 0, 147 => 0, 148 => 0, 149 => 0, 150 => 0, 151 => 0, 152 => 0, 153 => 0, 154 => 0, 155 => 0, 156 => 0, 157 => 1, 158 => 1, 159 => 1, 160 => 0, 161 => 0, 
162 => 0, 163 => 0, 164 => 0, 165 => 0, 166 => 0, 167 => 0, 168 => 0, 169 => 0, 170 => 0, 171 => 0, 172 => 0, 173 => 0, 174 => 0, 175 => 0, 176 => 0, 177 => 0, 178 => 0, 179 => 0, 180 => 0, 181 => 0, 182 => 0, 183 => 0, 184 => 0, 185 => 0, 186 => 0, 187 => 0, 188 => 0, 189 => 0, 190 => 0, 191 => 0, 192 => 0, 193 => 1, 194 => 0, 195 => 0, 196 => 0, 197 => 0, 198 => 0, 199 => 0, 200 => 0, 201 => 0, 202 => 0, 203 => 0, 204 => 0, 205 => 0, 206 => 0, 207 => 0, 208 => 0, 209 => 0, 210 => 0, 211 => 0, 212 => 0, 213 => 0, 214 => 0, 215 => 0, 216 => 0, 217 => 0, 218 => 0, 219 => 0, 220 => 0, 221 => 0, 222 
=> 0, 223 => 0, 224 => 0, 225 => 0, 226 => 0, 227 => 1, 228 => 1, 229 => 1, 230 => 0, 231 => 0, 232 => 0, 233 => 0, 234 => 0, 235 => 0, 236 => 0, 237 => 0, 238 => 0, 239 => 0, 240 => 0, 241 => 0, 242 => 0, 243 => 0, 244 => 0, 245 => 0, 246 => 0, 247 => 0, 248 => 0, 249 => 0, 250 => 0, 251 => 0, 252 => 0, 253 => 0, 254 => 0, 255 => 0, 256 => 0, 257 => 0, 258 => 0, 259 => 0, 260 => 0, 261 => 0, 262 => 0, 263 => 1, 264 => 0, 265 => 0, 266 => 0, 267 => 
0, 268 => 0, 269 => 0, 270 => 0, 271 => 0, 272 => 0, 273 => 0, 274 => 0, 275 => 0, 276 => 0, 277 => 0, 278 => 0, 279 => 0, 280 => 0, 281 => 0, 282 => 0, 283 => 0, 284 => 0, 285 => 0, 286 => 0, 287 => 0, 288 => 0, 289 => 0, 290 => 0, 291 => 0, 292 => 0, 293 => 0, 294 => 0, 295 => 0, 296 => 1, 297 => 1, 298 => 1, 299 => 0, 300 => 0, 301 => 0, 302 => 0, 303 => 0, 304 => 0, 305 => 0, 306 => 0, 307 => 0, 308 => 0, 309 => 0, 310 => 1, 311 => 1, 312 => 1, 
313 => 1, 314 => 1, 315 => 1, 316 => 1, 317 => 1, 318 => 1, 319 => 1, 320 => 1, 321 => 1, 322 => 1, 323 => 0, 324 => 0, 325 => 0, 326 => 0, 327 => 0, 328 => 0, 329 => 0, 330 => 0, 331 => 0, 332 => 1, 333 => 1, 334 => 1, 335 => 0, 336 => 0, 337 => 0, 338 => 0, 339 => 0, 340 => 0, 341 => 0, 342 => 0, 343 => 0, 344 => 0, 345 => 0, 346 => 1, 347 => 1, 348 => 1, 349 => 1, 350 => 1, 351 => 1, 352 => 1, 353 => 1, 354 => 1, 355 => 1, 356 => 1, 357 => 1, 358 => 1, 359 => 0, 360 => 0, 361 => 0, 362 => 0, 363 => 0, 364 => 0, 365 => 0, 366 => 0, 367 => 0, 368 => 0, 369 => 0, 370 => 0, 371 => 1, 372 => 0, 373 
=> 0, 374 => 0, 375 => 0, 376 => 0, 377 => 0, 378 => 0, 379 => 0, 380 => 0, 381 => 0, 382 => 0, 383 => 0, 384 => 0, 385 => 0, 386 => 0, 387 => 0, 388 => 0, 389 => 0, 390 => 0, 391 => 0, 392 => 0, 393 => 0, 394 => 0, 395 => 0, 396 => 0, 397 => 0, 398 => 0, 399 => 0, 400 => 0, 401 => 0, 402 => 0, 403 => 0, 404 => 0, 405 => 0, 406 => 0, 407 => 1, 408 => 1, 409 => 1, 410 => 0, 411 => 0, 412 => 0, 413 => 0, 414 => 0, 415 => 0, 416 => 0, 417 => 0, 418 => 
0, 419 => 0, 420 => 0, 421 => 0, 422 => 0, 423 => 0, 424 => 0, 425 => 0, 426 => 0, 427 => 0, 428 => 0, 429 => 0, 430 => 0, 431 => 0, 432 => 0, 433 => 0, 434 => 0, 435 => 0, 436 => 0, 437 => 0, 438 => 0, 439 => 0, 440 => 0, 441 => 0, 442 => 0, 443 => 0, 444 => 0, 445 => 1, 446 => 0, 447 => 0, 448 => 0, 449 => 0, 450 => 0, 451 => 0, 452 => 0, 453 => 0, 454 => 0, 455 => 0, 456 => 0, 457 => 0, 458 => 0, 459 => 0, 460 => 0, 461 => 0, 462 => 0, 463 => 0, 
464 => 0, 465 => 0, 466 => 0, 467 => 0, 468 => 0, 469 => 0, 470 => 0, 471 => 0, 472 => 0, 473 => 0, 474 => 0, 475 => 0, 476 => 0, 477 => 0, 478 => 0, 479 => 0, 480 => 0, 481 => 1, 482 => 1, 483 => 1, 484 => 0, 485 => 0, 486 => 0, 487 => 0, 488 => 0, 489 => 0, 490 => 0, 491 => 0, 492 => 0, 493 => 0, 494 => 0, 495 => 0, 496 => 0, 497 => 0, 498 => 0, 499 => 0, 500 => 0, 501 => 0, 502 => 0, 503 => 0, 504 => 0, 505 => 0, 506 => 0, 507 => 0, 508 => 0, 509 => 0, 510 => 0, 511 => 0, 512 => 0, 513 => 0, 514 => 0, 515 => 0, 516 => 0, 517 => 1, 518 => 1, 519 => 1, 520 => 0, 521 => 0, 522 => 0, 523 => 0, 524 
=> 0, 525 => 0, 526 => 0, 527 => 0, 528 => 0, 529 => 0, 530 => 0, 531 => 0, 532 => 0, 533 => 0, 534 => 0, 535 => 0, 536 => 0, 537 => 0, 538 => 0, 539 => 0, 540 => 0, 541 => 0, 542 => 0, 543 => 0, 544 => 0, 545 => 0, 546 => 0, 547 => 0, 548 => 0, 549 => 0, 550 => 0, 551 => 0, 552 => 0, 553 => 0, 554 => 0, 555 => 1, 556 => 1, 557 => 1, 558 => 1, 559 => 0, 560 => 0, 561 => 0, 562 => 0, 563 => 0, 564 => 0, 565 => 0, 566 => 0, 567 => 0, 568 => 0, 569 => 
0, 570 => 0, 571 => 0, 572 => 0, 573 => 0, 574 => 0, 575 => 0, 576 => 0, 577 => 0, 578 => 0, 579 => 0, 580 => 0, 581 => 0, 582 => 0, 583 => 0, 584 => 0, 585 => 0, 586 => 0, 587 => 0, 588 => 0, 589 => 0, 590 => 0, 591 => 1, 592 => 1, 593 => 1, 594 => 1, 595 => 0, 596 => 0, 597 => 0, 598 => 0, 599 => 0, 600 => 0, 601 => 0, 602 => 0, 603 => 0, 604 => 0, 605 => 0, 606 => 0, 607 => 0, 608 => 0, 609 => 0, 610 => 0, 611 => 0, 612 => 0, 613 => 0, 614 => 0, 
615 => 0, 616 => 0, 617 => 0, 618 => 0, 619 => 0, 620 => 0, 621 => 0, 622 => 0, 623 => 0, 624 => 0, 625 => 0, 626 => 0, 627 => 0, 628 => 0, 629 => 0, 630 => 0, 631 => 0, 632 => 0, 633 => 0, 634 => 0, 635 => 0, 636 => 0, 637 => 0, 638 => 0, 639 => 0, 640 => 0, 641 => 0, 642 => 0, 643 => 0, 644 => 0, 645 => 0, 646 => 0, 647 => 0
);

constant rom_ball: rom_bitmap_ball := (
0 => 0, 1 => 0, 2 => 0, 3 => 0, 4 => 0, 5 => 0, 6 => 0, 7 => 1, 8 => 1, 9 => 1, 10 => 1, 11 => 1, 12 => 1, 13 => 0, 14 => 0, 15 => 0, 16 => 0, 17 => 0, 18 => 0, 19 => 0, 20 => 0, 21 => 0, 22 => 0, 23 => 0, 24 => 0, 25 => 1, 26 => 1, 27 => 1, 28 => 1, 29 => 1, 30 => 1, 31 => 1, 32 => 1, 33 => 1, 34 => 
1, 35 => 0, 36 => 0, 37 => 0, 38 => 0, 39 => 0, 40 => 0, 41 => 0, 42 => 0, 43 => 0, 44 => 1, 45 => 1, 46 => 1, 47 => 1, 48 => 1, 49 => 1, 50 => 1, 51 => 1, 52 => 1, 53 => 1, 54 => 1, 55 => 1, 56 => 0, 57 => 0, 58 => 0, 59 => 0, 60 => 0, 61 => 0, 62 => 0, 63 => 1, 64 => 1, 65 => 1, 66 => 1, 67 => 1, 68 => 1, 69 => 1, 70 => 1, 71 => 1, 72 => 1, 73 => 1, 74 => 1, 75 => 1, 76 => 1, 77 => 0, 78 => 0, 79 => 0, 80 => 0, 81 => 0, 82 => 1, 83 => 1, 84 => 1, 
85 => 1, 86 => 1, 87 => 1, 88 => 1, 89 => 1, 90 => 1, 91 => 1, 92 => 1, 93 => 1, 94 => 1, 95 => 1, 96 => 1, 97 => 1, 98 => 0, 99 => 0, 100 => 0, 101 => 1, 102 => 1, 103 => 1, 104 => 1, 105 => 1, 106 => 1, 107 => 1, 108 => 1, 109 => 1, 110 => 1, 111 => 1, 112 => 1, 113 => 1, 114 => 1, 115 => 1, 116 => 
1, 117 => 1, 118 => 1, 119 => 0, 120 => 0, 121 => 1, 122 => 1, 123 => 1, 124 => 1, 125 => 1, 126 => 1, 127 => 1, 128 => 1, 129 => 1, 130 => 1, 131 => 1, 132 => 1, 133 => 1, 134 => 1, 135 => 1, 136 => 1, 137 => 1, 138 => 1, 139 => 0, 140 => 1, 141 => 1, 142 => 1, 143 => 1, 144 => 1, 145 => 1, 146 => 1, 147 => 1, 148 => 1, 149 => 1, 150 => 1, 151 => 1, 152 => 1, 153 => 1, 154 => 1, 155 => 1, 156 => 1, 157 => 1, 158 => 1, 159 => 1, 160 => 1, 161 => 1, 
162 => 1, 163 => 1, 164 => 1, 165 => 1, 166 => 1, 167 => 1, 168 => 1, 169 => 1, 170 => 1, 171 => 1, 172 => 1, 173 => 1, 174 => 1, 175 => 1, 176 => 1, 177 => 1, 178 => 1, 179 => 1, 180 => 1, 181 => 1, 182 => 1, 183 => 1, 184 => 1, 185 => 1, 186 => 1, 187 => 1, 188 => 1, 189 => 1, 190 => 1, 191 => 1, 192 => 1, 193 => 1, 194 => 1, 195 => 1, 196 => 1, 197 => 1, 198 => 1, 199 => 1, 200 => 1, 201 => 1, 202 => 1, 203 => 1, 204 => 1, 205 => 1, 206 => 1, 207 => 1, 208 => 1, 209 => 1, 210 => 1, 211 => 1, 212 => 1, 213 => 1, 214 => 1, 215 => 1, 216 => 1, 217 => 1, 218 => 1, 219 => 1, 220 => 1, 221 => 1, 222 
=> 1, 223 => 1, 224 => 1, 225 => 1, 226 => 1, 227 => 1, 228 => 1, 229 => 1, 230 => 1, 231 => 1, 232 => 1, 233 => 1, 234 => 1, 235 => 1, 236 => 1, 237 => 1, 238 => 1, 239 => 1, 240 => 1, 241 => 1, 242 => 1, 243 => 1, 244 => 1, 245 => 1, 246 => 1, 247 => 1, 248 => 1, 249 => 1, 250 => 1, 251 => 1, 252 => 1, 253 => 1, 254 => 1, 255 => 1, 256 => 1, 257 => 1, 258 => 1, 259 => 1, 260 => 0, 261 => 1, 262 => 1, 263 => 1, 264 => 1, 265 => 1, 266 => 1, 267 => 
1, 268 => 1, 269 => 1, 270 => 1, 271 => 1, 272 => 1, 273 => 1, 274 => 1, 275 => 1, 276 => 1, 277 => 1, 278 => 1, 279 => 0, 280 => 0, 281 => 1, 282 => 1, 283 => 1, 284 => 1, 285 => 1, 286 => 1, 287 => 1, 288 => 1, 289 => 1, 290 => 1, 291 => 1, 292 => 1, 293 => 1, 294 => 1, 295 => 1, 296 => 1, 297 => 1, 298 => 1, 299 => 0, 300 => 0, 301 => 0, 302 => 1, 303 => 1, 304 => 1, 305 => 1, 306 => 1, 307 => 1, 308 => 1, 309 => 1, 310 => 1, 311 => 1, 312 => 1, 
313 => 1, 314 => 1, 315 => 1, 316 => 1, 317 => 1, 318 => 0, 319 => 0, 320 => 0, 321 => 0, 322 => 0, 323 => 1, 324 => 1, 325 => 1, 326 => 1, 327 => 1, 328 => 1, 329 => 1, 330 => 1, 331 => 1, 332 => 1, 333 => 1, 334 => 1, 335 => 1, 336 => 1, 337 => 0, 338 => 0, 339 => 0, 340 => 0, 341 => 0, 342 => 0, 343 => 0, 344 => 1, 345 => 1, 346 => 1, 347 => 1, 348 => 1, 349 => 1, 350 => 1, 351 => 1, 352 => 1, 353 => 1, 354 => 1, 355 => 1, 356 => 0, 357 => 0, 358 => 0, 359 => 0, 360 => 0, 361 => 0, 362 => 0, 363 => 0, 364 => 0, 365 => 1, 366 => 1, 367 => 1, 368 => 1, 369 => 1, 370 => 1, 371 => 1, 372 => 1, 373 
=> 1, 374 => 1, 375 => 0, 376 => 0, 377 => 0, 378 => 0, 379 => 0, 380 => 0, 381 => 0, 382 => 0, 383 => 0, 384 => 0, 385 => 0, 386 => 0, 387 => 1, 388 => 1, 389 => 1, 390 => 1, 391 => 1, 392 => 1, 393 => 0, 394 => 0, 395 => 0, 396 => 0, 397 => 0, 398 => 0, 399 => 0
);
		function to_std_logic(i : integer) return std_logic is
	begin
		 if i = 0 then
			  return '0';
		 end if;
		 return '1';
	end function;
	
	constant H_ACTIVE_AREA: integer := 800;	
	constant H_END_FP: integer := 856;--FP - FRONT PORCH	
	constant H_END_SPULSE: integer := 976;--SYNC PULSE
	constant H_END_BP: integer := 1040;-- BACK PORCH
	
	--same as above, but for vertical area
	constant V_ACTIVE_AREA: integer := 600;	
	constant V_END_FP: integer := 637;--FP - FRONT PORCH	
	constant V_END_SPULSE: integer := 643;
	constant V_END_BP: integer := 666;
	
	--constants for paddle and ball size
	constant P_HEIGHT: integer := 140;
	constant P_WIDTH: integer := 15;
	constant B_RADIUS: integer := 10; --16 PER SIDE
	constant N_WIDTH: integer := 2;
	constant N_HEIGHT: integer := 20;
	constant N_GAP:	 integer := 10;
	
	constant SCORE_X: integer := H_ACTIVE_AREA/4;
	constant SCORE_Y: integer := V_ACTIVE_AREA/4;
	constant TILE: integer := 12;
	constant GAP: integer := 3;
	constant SCORE_WIDTH: integer := TILE*6 + 2*GAP;
	constant SCORE_HEIGHT: integer:= TILE*4 + GAP;

	constant TITLE_WIDTH: integer := 200;
	constant TITLE_HEIGHT: integer := 45;
	constant TITLE_GAP_X: integer := 36;
	constant PONG_WIDTH: integer := 198;
	
	constant OPTION_WIDTH: integer := 164;
	constant OPTION_HEIGHT: integer := 18;--constant ARROW_HEIGHT: integer:= 18;
	
	constant ARROW_WIDTH: integer := 36;
	
	constant TITLE_X: integer := H_ACTIVE_AREA/2 - TITLE_WIDTH/2 - PONG_WIDTH/2 - TITLE_GAP_X/2;
	constant TITLE_Y: integer := V_ACTIVE_AREA/4;
	constant TITLE_GAP: integer := TITLE_Y;
	constant OPTION_GAP:		integer := 20;
	constant OPTION_X: integer := H_ACTIVE_AREA/2 - OPTION_WIDTH/2; 
	constant OPTION_Y: integer:= TITLE_Y + TITLE_HEIGHT + TITLE_GAP;
	
	constant OPTION_LIMIT: integer := 2951;--3599;2
	constant TITLE_LIMIT: integer := 8999;
	constant TITLE_PONG: integer 	:= 8909;
	constant ARROW_LIMIT: integer := 647;
	
	constant BORDER_WIDTH: integer := 5;
	
	constant JS1_DELAY: integer := 1666500;--1250000;--25ms (40ms 40upd/s) --2500000; --50ms(20 upd/s) 
		
	--counts to keep track of position of the actual pixel being rended
	signal r_count_x: integer := 0;	--hs 
	signal r_count_y: integer := 0;	--vs
	
	--vector representation from the above counter
	signal v_count_y: std_logic_vector(9 downto 0);
	
	--pulses for HS and VS drive signals to proper show image
	signal w_HS: std_logic;	
	signal w_VS: std_logic;
	
	--hints for active pixels on the display
	signal w_HD_active: std_logic;	
	signal w_VD_active: std_logic;
	--for control draw
	signal w_draw_paddle1: std_logic := '0';	
	signal w_draw_paddle2: std_logic := '0';	
	signal w_draw_ball: std_logic := '0';
	signal w_draw_border: std_logic := '0';	
	signal w_draw_net: std_logic := '0';
	
	signal w_ball_x: integer range 0 to H_ACTIVE_AREA := H_ACTIVE_AREA/2;
	signal w_ball_Y: integer range 0 to V_ACTIVE_AREA := V_ACTIVE_AREA/2;
	--signal ball_count: integer := 0;

	signal w_render: std_logic;
	signal w_inBall: std_logic;	
	signal w_inBorder: std_logic;	
	signal w_inPaddle1: std_logic;	
	signal w_inPaddle2: std_logic;
	signal w_inNet: std_logic;	
	signal w_inDisplay: std_logic;
	--for menu
	signal w_inTitle: std_logic 	:= '0';	
	signal w_inPong: std_logic 	:= '0';
	signal w_inOption1: std_logic := '0';	
	signal w_inOption2: std_logic := '0';	
	signal w_arrow_in_option2: std_logic := '0';
	signal w_arrow_in_option1: std_logic := '0';
	
	signal option1_count: integer :=0;
	signal option2_count: integer :=0;
	signal title_count: integer := 0;	
	signal pong_count: integer := 0;	
	signal arrow_count: integer := 0;
	
	signal w_draw_arrow: std_logic := '0';
	signal w_draw_title: std_logic := '0';	
	signal w_draw_pong: std_logic := '0';
	signal w_draw_option1: std_logic := '0';
	signal w_draw_option2: std_logic := '0';
	
	signal 	w_paddle1_y: integer range 0 to V_ACTIVE_AREA - P_HEIGHT := V_ACTIVE_AREA/2 - P_HEIGHT/2;
	constant w_paddle1_x: integer := 5 + BORDER_WIDTH;
	signal 	w_paddle2_y: integer range 0 to V_ACTIVE_AREA - P_HEIGHT := V_ACTIVE_AREA/2 - P_HEIGHT/2;
	constant w_paddle2_x: integer := H_ACTIVE_AREA - P_WIDTH - w_paddle1_x;
	
	constant w_ball_vel_x:	integer range 0 to 10 := 5;		
	constant w_ball_vel_y:	integer range 0 to 10 := 5;
	signal w_vel_dir_x: std_logic := '1';	
	signal w_vel_dir_y: std_logic := '1';	
	-- for 4-point collision detection
	signal w_collision_in_left: std_logic;	
	signal w_collision_in_right: std_logic;
	signal w_collision_in_both_x: std_logic;
	
	signal w_collision_in_top: std_logic;	
	signal w_collision_in_bottom: std_logic;
	signal w_collision_in_both_y: std_logic;
	
	signal collide_in_left: std_logic;
	signal collide_in_right: std_logic;
	signal collide_in_top: std_logic;
	signal collide_in_bottom: std_logic;
	signal w_collide_in_p1: std_logic := '0';
	signal w_collide_in_p2: std_logic := '0';	
	signal w_collide_mid_to_bottom: std_logic := '0';
	signal w_collide_mid_to_top: std_logic := '0';
	signal w_collide_mid_to_bottom_p2: std_logic := '0';
	signal w_collide_mid_to_top_p2: std_logic := '0';
	
	signal w_reset_collision: std_logic;
	signal w_is_drawing: std_logic;
	signal w_one_per_frame: std_logic := '0';	
	
	signal w_joystick_p1: integer range 0 to 64 := 31;--middle or 0	
	signal w_js1_UP: std_logic;
	signal w_js1_DOWN: std_logic;
	
	signal w_joystick_p2: integer range 0 to 64 := 31;--middle or 0	
	signal w_js2_UP: std_logic;
	signal w_js2_DOWN: std_logic;
	
	signal w_in_range: std_logic;
	signal w_js1_count: integer := 0;
	signal w_versus_com: std_logic;
	signal w_in_range_p2: std_logic;
	signal w_js2_count: integer := 0;
	signal w_increment: integer := 0;
	
	signal w_do_wall_sound : std_logic := '0' ;	
	signal w_do_paddle_sound : std_logic := '0' ;
	signal w_do_point_sound : std_logic := '0' ;	
	signal w_do_select_sound : std_logic := '0' ;
	
	signal w_render_active: std_logic := '0';
	signal w_default_option: std_logic := '0';
	signal w_draw_menu:		std_logic := '0';
	signal w_select: std_logic := '0';
	signal w_score_p1 : integer := 0;	
	signal w_score_p2 : integer := 0;
	signal w_draw_score_p1: std_logic := '0';
	signal w_draw_score_p2: std_logic := '0';
	signal w_active_score: std_logic := '0';
	
	--signal w_delay_play: integer := 0;

	type t_game is (s_menu, s_play);
	
	signal game_flow: t_game := s_menu;
begin

	--for joystick
	w_joystick_p1 <= to_integer(unsigned(i_joystick_p1));
	w_js1_UP <= '1' when w_joystick_p1 > 36 else '0';	
	w_js1_DOWN <= '1' when w_joystick_p1 < 27 else '0';
	w_in_range <= '1' when w_paddle1_y > BORDER_WIDTH and w_paddle1_y < V_ACTIVE_AREA - P_HEIGHT - BORDER_WIDTH else '0';
	--paddle2
	w_joystick_p2 <= to_integer(unsigned(i_joystick_p2));
	w_js2_DOWN <= '1' when w_joystick_p2 > 36 else '0';	
	w_js2_UP <= '1' when w_joystick_p2 < 27 else '0';
	w_in_range_p2 <= '1' when w_paddle2_y >= BORDER_WIDTH and w_paddle2_y <= V_ACTIVE_AREA - P_HEIGHT - BORDER_WIDTH  else '0';
	
	--for draw
	v_count_y <= std_logic_vector(to_unsigned(r_count_y, v_count_y'length));	
	w_inBorder <= '1' when (r_count_x >= 0  and r_count_x <= BORDER_WIDTH) or (r_count_x >= H_ACTIVE_AREA - BORDER_WIDTH and r_count_x <= H_ACTIVE_AREA) or 
	(r_count_y >= 0 and r_count_y <= BORDER_WIDTH) or (r_count_y >= V_ACTIVE_AREA - BORDER_WIDTH and r_count_y <= V_ACTIVE_AREA) else '0';									  
	w_inBall <= '1' when r_count_x >= w_ball_x - B_RADIUS and r_count_x <= w_ball_x + B_RADIUS  -- left and right side, respectively
	and r_count_y >= w_ball_y - B_RADIUS and r_count_y <= w_ball_y + B_RADIUS -- top and bottom side , //
	else '0';
	w_inPaddle1 <= '1' when r_count_x >= w_paddle1_x and r_count_x <= w_paddle1_x + P_WIDTH and 
									r_count_y >= w_paddle1_y and r_count_y <= w_paddle1_y + P_HEIGHT else '0';
	w_inPaddle2 <= '1' when r_count_x >= w_paddle2_x and r_count_x <= w_paddle2_x + P_WIDTH and 
									r_count_y >= w_paddle2_y and r_count_y <= w_paddle2_y + P_HEIGHT else '0';								
	w_inNet <= '1' when (v_count_y(4) = '0' and (r_count_x >= H_ACTIVE_AREA/2 - N_WIDTH/2 and 
															  r_count_x <= H_ACTIVE_AREA/2 + N_WIDTH/2) ) else '0';
	
	-- ball collision
	w_is_drawing <= '1' when (w_draw_border = '1') or (w_draw_paddle1 = '1') or (w_draw_paddle2 = '1') else '0';
	collide_in_left <= '1' when w_is_drawing = '1' and r_count_x = w_ball_x - B_RADIUS and r_count_y = w_ball_y else '0';
	collide_in_right <= '1' when w_is_drawing = '1' and (r_count_x = w_ball_x + B_RADIUS and r_count_y = w_ball_y) else '0';												
	collide_in_top <= '1' when w_is_drawing = '1' and r_count_x = w_ball_x and r_count_y = w_ball_y - B_RADIUS else '0';											
	collide_in_bottom <= '1' when w_is_drawing = '1' and r_count_x = w_ball_x and r_count_y = w_ball_y + B_RADIUS else '0';	
	w_collision_in_both_x <= '1' when w_collision_in_left = '1' and w_collision_in_right = '1' else '0';
	w_collision_in_both_y <= '1' when w_collision_in_bottom = '1' and w_collision_in_top = '1' else '0';
	
	--paddle collision
	w_collide_in_p1 <= '1' when w_ball_x - B_RADIUS <= w_paddle1_x + P_WIDTH  else '0';	
	w_collide_in_p2 <= '1' when w_ball_x + B_RADIUS >= w_paddle2_x else '0';
	w_collide_mid_to_bottom <= '1' when (w_ball_y >= w_paddle1_y + P_HEIGHT/2 and w_ball_y < w_paddle1_y + P_HEIGHT) else '0';-- '1' -> (middle to bottom)
	w_collide_mid_to_top <= '1' when (w_ball_y >= w_paddle1_y and w_ball_y < w_paddle1_y + P_HEIGHT/2) else '0';-- 
	w_collide_mid_to_bottom_p2 <= '1' when (w_ball_y >= w_paddle2_y + P_HEIGHT/2 and w_ball_y < w_paddle2_y + P_HEIGHT) else '0';-- '1' -> (middle to bottom)
	w_collide_mid_to_top_p2 <= '1' when (w_ball_y >= w_paddle2_y and w_ball_y < w_paddle2_y + P_HEIGHT/2) else '0';
	
	--for menu--								 
	w_inPong <= '1' when r_count_x > TITLE_X and r_count_x <= TITLE_X + PONG_WIDTH and
								r_count_y > TITLE_Y and r_count_y <= TITLE_Y + TITLE_HEIGHT else '0';
	
	w_inTitle <= '1' when r_count_x > TITLE_X + PONG_WIDTH + TITLE_GAP_X and 
								 r_count_x <= TITLE_X + PONG_WIDTH + TITLE_GAP_X + TITLE_WIDTH and
								 r_count_y > TITLE_Y and r_count_y <= TITLE_Y + TITLE_HEIGHT else '0';
	
	w_inOption1 <= '1' when r_count_x > OPTION_X and r_count_x <= OPTION_X + OPTION_WIDTH and
									r_count_y >= OPTION_Y and r_count_y <= OPTION_Y + OPTION_HEIGHT else '0';
									
	w_arrow_in_option1 <= '1' when r_count_x > OPTION_X + OPTION_WIDTH and 
											 r_count_x <= OPTION_X + OPTION_WIDTH + ARROW_WIDTH and
											 r_count_y > OPTION_Y and r_count_y <= OPTION_Y + OPTION_HEIGHT else '0';
	
	w_inOption2 <= '1' when r_count_x > OPTION_X and r_count_x <= OPTION_X + OPTION_WIDTH and
									r_count_Y > OPTION_Y + OPTION_HEIGHT*2 and r_count_y <= OPTION_Y + OPTION_HEIGHT*3 else '0';    
									
	w_arrow_in_option2 <= '1' when r_count_x > OPTION_X + OPTION_WIDTH and 
											 r_count_x <= OPTION_X + OPTION_WIDTH + ARROW_WIDTH and
											 r_count_y >= OPTION_Y + OPTION_HEIGHT*2 
										and r_count_y <= OPTION_Y + OPTION_HEIGHT*3 else '0';
	
	process(i_clk)
	begin
		if rising_edge(i_clk) then
			case game_flow is 
				when s_menu =>
					w_active_score <= '0';
					w_score_p1 <= 0;
					w_score_p2 <= 0;	
					w_draw_border <= '0';
					w_draw_paddle1 <= '0';
					w_draw_paddle2 <= '0';
					w_draw_net <= '0';
					w_draw_ball <= '0';
					w_do_point_sound <= '0';
					if w_js1_UP = '1' then
						w_default_option <= '0';
					elsif w_js1_DOWN = '1' then
						w_default_option <= '1'; 
					end if;
					--one player, vs computer
					if w_select = '1' and w_default_option = '0' then
						game_flow <= s_play;
						w_versus_com <= '1';
						w_do_select_sound <= '1';
					elsif w_select = '1' and w_default_option = '1' then
						game_flow <= s_play;
						w_versus_com <= '0';
						w_do_select_sound <= '1';
					end if;
					
					--for draw menu
					if r_count_y = V_ACTIVE_AREA - 1 and r_count_x = H_ACTIVE_AREA -1 then
						pong_count <= 0;
					else
						if w_inPong = '1' and pong_count <= TITLE_PONG then
							pong_count <= pong_count + 1;
							w_draw_pong <= to_std_logic(rom_pong(pong_count));
						else
							w_draw_pong <= '0';
						end if;
					end if;
					
					if r_count_y = V_ACTIVE_AREA - 1 and r_count_x = H_ACTIVE_AREA -1 then
						title_count <= 0;
					else
						if w_inTitle = '1' and title_count <= TITLE_LIMIT then
							title_count <= title_count + 1;
							w_draw_title <= to_std_logic(rom_game(title_count));
						else
							w_draw_title <= '0';
						end if;
					end if;
						
					if r_count_y = V_ACTIVE_AREA - 1 and r_count_x = H_ACTIVE_AREA -1 then
						option1_count <= 0;
					else
						if w_inOption1 = '1' and option1_count <= OPTION_LIMIT then
							option1_count <= option1_count + 1;
							w_draw_option1 <= to_std_logic(rom_option_1(option1_count));
						else
							w_draw_option1 <= '0';
						end if;
					end if;	
					
					if r_count_y = V_ACTIVE_AREA - 1 and r_count_x = H_ACTIVE_AREA -1 then
						option2_count <= 0;
					else
						if w_inOption2 = '1' and option2_count <= OPTION_LIMIT then
							option2_count <= option2_count + 1;
							w_draw_option2 <= to_std_logic(rom_option_2(option2_count));
						else
							w_draw_option2 <= '0';
						end if;
					end if;
					
					if r_count_y = V_ACTIVE_AREA - 1 and r_count_x = H_ACTIVE_AREA -1 then
						arrow_count <= 0;
					else
						if w_default_option = '1' then
							
							if w_arrow_in_option2 = '1' and arrow_count <= ARROW_LIMIT then
								arrow_count <= arrow_count + 1;
								w_draw_arrow <= to_std_logic(rom_arrow(arrow_count));
							else
								w_draw_arrow <= '0';
							end if;
						else
							if w_arrow_in_option1 = '1' and arrow_count <= ARROW_LIMIT then
								arrow_count <= arrow_count + 1;
								w_draw_arrow <= to_std_logic(rom_arrow(arrow_count));
							else
								w_draw_arrow <= '0';
							end if;
						end if;
					end if;
					
				
				when s_play =>
					w_do_select_sound <= '0';
					w_active_score <= '1';
					
					if w_inBorder = '1' then
						w_draw_border <= '1';
					else 
						w_draw_border <= '0';
					end if;
					
					if w_inPaddle1 = '1' then
						w_draw_paddle1 <= '1';
					else
						w_draw_paddle1 <= '0';
					end if;
				
					if w_inPaddle2 = '1' then
						w_draw_paddle2 <= '1';
					else
						w_draw_paddle2 <= '0';
					end if;
					
					if w_inNet = '1' then
						w_draw_net <= '1';
					else 
						w_draw_net <= '0';
					end if;
					
					if w_inBall = '1' then
						w_draw_ball <= '1';
					else
						w_draw_ball <= '0';
					end if;
					--end draw section
					
					if w_js1_count < JS1_DELAY then
						w_js1_count <= w_js1_count + 1;
					else
						w_js1_count <= 0;
						
						if w_in_range = '1' then
							if w_js1_UP = '1' then
							 w_paddle1_y <= w_paddle1_y - 10;
							elsif w_js1_DOWN = '1' then
							 w_paddle1_y <= w_paddle1_y + 10;
							end if;
						elsif w_paddle1_y <= BORDER_WIDTH and w_js1_DOWN = '1' then
							w_paddle1_y <= w_paddle1_y + 10;
						elsif w_paddle1_y >= V_ACTIVE_AREA - P_HEIGHT  - BORDER_WIDTH and w_js1_UP = '1' then
							w_paddle1_y <= w_paddle1_y - 10;
						end if;
					end if;
					
					if w_js2_count < JS1_DELAY then
						w_js2_count <= w_js2_count + 1;
					else
						w_js2_count <= 0;
							if w_versus_com = '1' then
								if i_difficulty = "00" then
									w_increment <= (w_ball_y - (w_paddle2_y + P_HEIGHT/2))/8;
								elsif i_difficulty = "01" then
									w_increment <= (w_ball_y - (w_paddle2_y + P_HEIGHT/2))/4;
								elsif i_difficulty = "10" then  
									w_increment <= (w_ball_y - (w_paddle2_y + P_HEIGHT/2))/2;
								else
									w_increment <= (w_ball_y - (w_paddle2_y + P_HEIGHT/2))/8;
								end if;
								if w_in_range_p2 = '1' then
									w_paddle2_y <= w_paddle2_y + w_increment;
								elsif w_paddle2_y <= BORDER_WIDTH and w_increment > 0 then
									w_paddle2_y <= w_paddle2_y + w_increment;
								elsif w_paddle2_y >= V_ACTIVE_AREA - P_HEIGHT - BORDER_WIDTH and w_increment < 0 then
									w_paddle2_y <= w_paddle2_y + w_increment;
								end if;
							else
								if w_in_range_p2 = '1' then
									if w_js2_UP = '1' then
									 w_paddle2_y <= w_paddle2_y - 10;
									elsif w_js2_DOWN = '1' then
									 w_paddle2_y <= w_paddle2_y + 10;
									end if;
								elsif w_paddle2_y <= BORDER_WIDTH and w_js2_DOWN = '1' then
									w_paddle2_y <= w_paddle2_y + 10;
								elsif w_paddle2_y >= V_ACTIVE_AREA - P_HEIGHT - BORDER_WIDTH and w_js2_UP = '1' then
									w_paddle2_y <= w_paddle2_y - 10;
								end if;
							end if;
					end if;
					
					if w_reset_collision = '1' then
						w_collision_in_left <= '0';				
						w_collision_in_right <= '0';
						w_collision_in_top <= '0';
						w_collision_in_bottom <= '0';
					else 
					
						if collide_in_left = '1' then
							w_collision_in_left <= '1';
						end if;
						
						if collide_in_right = '1' then
							w_collision_in_right <= '1';
						end if;
						
						if collide_in_top = '1' then
							w_collision_in_top <= '1';
						end if;
						
						if collide_in_bottom = '1' then
							w_collision_in_bottom <= '1';
						end if;
						
					end if;
					
					if (r_count_y /= V_ACTIVE_AREA - 1) OR (r_count_x /= H_ACTIVE_AREA - 1) then
						w_reset_collision <= '0';
						if w_one_per_frame = '0' then
							w_one_per_frame <= '1';
							if w_collision_in_both_x = '0' then
								--'1' -> go to left, '0' -> go to right
								if w_vel_dir_x = '1' then
									w_ball_x <= w_ball_x - w_ball_vel_x;
								else
									w_ball_x <= w_ball_x + w_ball_vel_x;
								end if;
								
								if w_collision_in_left = '1' then
									--go to right
									w_vel_dir_x <= '0';
									
									if w_collide_mid_to_bottom = '1' and w_collide_in_p1 = '1' then
										--go to right and bottom
										w_vel_dir_y <= '0';
										w_do_paddle_sound <= '1';
									elsif w_collide_in_p1 = '1' and w_collide_mid_to_top = '1' then
										--go to right and top
										w_vel_dir_y <= '1';
										w_do_paddle_sound <= '1';
									end if;
								elsif w_collision_in_right = '1' then 
									--go to left
									w_vel_dir_x <= '1';
									
									if w_collide_mid_to_bottom_p2 = '1' and w_collide_in_p2 = '1' then
										--go to left and bottom
										w_vel_dir_y <= '0';
										w_do_paddle_sound <= '1';
									elsif w_collide_in_p2 = '1' and w_collide_mid_to_top_p2 = '1' then
										--go to right and top
										w_vel_dir_y <= '1';
										w_do_paddle_sound <= '1';
									end if;
								else
									w_do_paddle_sound <= '0';
								end if;
							
							end if;
							
							if w_collision_in_both_y = '0' then
								--'1' -> up , 0' -> down
								if w_vel_dir_y = '1' then
									w_ball_y <= w_ball_y - w_ball_vel_y;
								else 
									w_ball_y <= w_ball_y + w_ball_vel_y;
								end if;
								
								if w_collision_in_top = '1' then
									--go to down
									w_vel_dir_y <= '0';
									w_do_wall_sound <= '1';
								elsif w_collision_in_bottom = '1' then
									--go up to
									w_vel_dir_y <= '1';
									w_do_wall_sound <= '1';
								else
									w_do_wall_sound <= '0';
								end if;
							end if;
								
							if w_ball_x - B_RADIUS <= BORDER_WIDTH then --collide in border of ps1 then point for ps2
								w_ball_x <= H_ACTIVE_AREA/2;
								w_ball_y <= V_ACTIVE_AREA/2;
		--						w_vel_dir_x <= '0';
								w_do_point_sound <= '1';
								w_score_p2 <= w_score_p2 + 1;
							elsif w_ball_x + B_RADIUS >= H_ACTIVE_AREA - BORDER_WIDTH then 
								w_ball_x <= H_ACTIVE_AREA/2;
								w_ball_y <= V_ACTIVE_AREA/2;
								w_vel_dir_x <= '1';
								w_do_point_sound <= '1';
								w_score_p1 <= w_score_p1 + 1;
								--score fot ps1
							else 
								w_do_point_sound <= '0';
							end if;
		--					
						end if;
						
						if w_score_p2 = 10 or w_score_p1 = 10 then
							game_flow <= s_menu;
						end if;
					else
						w_reset_collision <= '1';
						w_one_per_frame <= '0';							
					end if;
				
				when others => game_flow <= s_menu;	
			end case;
		end if;	
	end process;
	
	debounce: entity work.Debounce_Switch
	port map(
		i_Clk 	=> i_clk,
		i_Switch => i_select,
		o_Switch => w_select
	);
	
	--VGA
	w_render <= '1' when (w_draw_ball = '1') or (w_draw_border = '1') or 
								(w_draw_paddle1 = '1') or (w_draw_paddle2 = '1') or
								(w_draw_net = '1') or (w_draw_menu = '1') OR
								(w_draw_arrow = '1') or (w_draw_option1 = '1') or
								(w_draw_option2 = '1') or (w_draw_score_p1 = '1') or 
								(w_draw_score_p2 = '1') or (w_draw_title = '1') or 
								(w_draw_pong = '1') else '0';
								
	w_inDisplay <= '1' when w_HD_active = '1' and w_VD_active = '1' else '0';

	o_R0 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_R1 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_R2 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_G0 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_G1 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_G2 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_B0 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	o_B1 <= '1' when w_inDisplay = '1' and w_render = '1' else '0';
	
	o_HS <= w_HS;	
	o_VS <= w_VS;
	
	vga_controller: entity work.vga_controller
	generic map(
		--FREQLIMIT: integer;
		H_ACTIVE_AREA => H_ACTIVE_AREA,
		H_END_FP			=> H_END_FP,
		H_END_SPULSE	=> H_END_SPULSE,
		H_END_BP			=> H_END_BP,
		V_ACTIVE_AREA	=> V_ACTIVE_AREA,
		V_END_FP			=> V_END_FP,
		V_END_SPULSE	=> V_END_SPULSE,
		V_END_BP			=> V_END_BP
	)
	port map(
		i_clk       => i_clk, 
		o_HS  		=> w_HS,
		o_VS			=> W_VS,
		o_HD_active	=> w_HD_active,
		o_VD_active => w_VD_active,
		o_col_count => r_count_x,
		o_row_count => r_count_y
	);
	
	p1_score: entity work.score_counter
	generic map(
		SCORE_X			=> SCORE_X,
		SCORE_Y			=> SCORE_Y,
		TILE				=>	TILE,
		GAP				=> GAP,
		SCORE_WIDTH		=> SCORE_WIDTH,
		SCORE_HEIGHT 	=>	SCORE_HEIGHT
	)
	port map(
		i_clk					=> i_clk,
		r_count_x   		=> r_count_x,
		r_count_y   		=> r_count_y,
		i_score     		=> w_score_p1,
		i_active_render	=> w_active_score,
		o_segment   		=> w_draw_score_p1
	);
	
	p2_score: entity work.score_counter
	generic map(
		SCORE_X 			=> H_ACTIVE_AREA/2 + H_ACTIVE_AREA/4  - SCORE_WIDTH,
		SCORE_Y			=> SCORE_Y,
		TILE				=>	TILE,
		GAP				=> GAP,
		SCORE_WIDTH		=> SCORE_WIDTH,
		SCORE_HEIGHT	=> SCORE_HEIGHT
	)
	port map(
		i_clk					=> i_clk,
		r_count_x   		=> r_count_x,
		r_count_y   		=> r_count_y,
		i_score     		=> w_score_p2,
		i_active_render	=> w_active_score,
		o_segment   		=> w_draw_score_p2
	);
	
	pong_sounds: entity work.sound_for_pong
	port map(
		i_clk 					=> i_clk,
		paddle_sound_collide => o_paddle_sound_collide,
		do_wall_sound			=> w_do_wall_sound,
		do_paddle_sound		=> w_do_paddle_sound,
		do_point_sound			=> w_do_point_sound,
		do_select_sound		=> w_do_select_sound
	);
	
end Behavioral;


